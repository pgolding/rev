BZh91AY&SY�)� l߀Py��g߰?���P�u  	"I�#F��4M44 �@h��h9�&L�0�&&��!�0# ����4�T��I��  4�i��&�&	��0`��"��L!=T���T�Sjz��  Q�0��1YT	b��Ň���	�
��bI�P����*����/H��]T$�Sub��M]eeEjP7{췚���2ZL&5`�\N�A,
�37�VRU�Ē4���<?�e�rc�L�?ܜ��b\�F\ W�`3��� q���c�I{c(U��w�YT"�J&�&di�𴶅ܔ[Ak��4��6�l�����0h��aЩu��*���j���W��,��0�$+J����ȦE�`օγjL���kd�%BR����&[�馆h̭8>��+��*Q)�fT����1]%�ť5 a��J��su!�-[� ��"l|��S~���P�G�8�&$˄����1 �q��[ģ��ܴ�ܡED��y�6��M�S]`)�FD�*u%��B�MJ��=;�R�K"t:���1�����=L��~��%��v�v����zu��J_)����pfń�MC]�O��`�,']O�Ǚ	�8��<����MX�3�ӢV�H���r�����(;Q`��2	~��R��\N�a�	���iD���t	L;�s����_�@ƺ�|0|��$�����'m���dT's���������ڹbl��D��А���ԯ��K@�M�u,��3�1xƫ��~�����APW9[vf��C��r��*|���,�-۷/�;���A�)����8<Y�F�aMWa��" �y�nV���H�
�1 �