BZh91AY&SY����R߀rpg���>� ?���a��                                           ;�@�EUJ��AUR�
�U*J�JB�U" B���UB$R��IU*�$��R�"RT��	J��IT)PJs�B� =����H�$P���D�x'�8C `���<�H������������n���
��#�     ��}�TxY��*��T�)�R�ggxm*��ܫ�4�Z�8Myj�S��U*�y�R�ۧ�Ԫ��Tx�W��W���T��   �BDJP��$I�/��I>�U�t�ڕ\f��ʽ�Ԫ�Y��*�<T����U��R��Rri^��x��Y�R���$����x��j���W�   wJ��R���۪�W���PW�J����ʧzܧ�UyjUsgy�U*�ފ�'z�Sy�J��W6U�n�W�^��W�   <�B��QP�����EB]歹]���5W-Uϻ���*�k��U]��U��UWv誩�Ϋ֪��I�qeUOniT�9�R����T��wU�   ��ʫl��U7�*�n�Us���P�Xs�Uw�UU�;��UW]�UAΪ���UT��%s������UO�   = UD�UJ��� ުU[�M�C���U�U+f��UR�9*�7U*�ۧmU9���j�۫�^��T;��RE#ê�i�V��_   4Χ����^Z�U댨*��UY��Z��K�}>��*���=ê���A��U[�O6���w��9W�UUɸ����   ��E%P�B�R�%T���"��w7<�U\m'{��ݺ��k��UJ�T�J��޳�Z���:�L�����q�US�ށR��U�O&��7K�   �����k�붼>�U{ʕݏg������o.��7|ܪx��*����S����|�χ����w��v��uK�              ?T�$����0�4ё��M&�)R��P�4�j �` 0�4?&�U  4     '�T�(�I        5?B�?*�Tѐa0@��&��%$��d�&�S�MM4=&F���b#�'�S�~g�~�އ���I�x��Ϟ�����z珕U@<�܏�U@>�����ETA� ����"���������u��_��?�������|��������������O�Ҩ��Q��/���I�ݓ�Ђ��x�����������z��ށET�g�=�V*�UR���b�p�e��Ēh��PS����1E��	���m�ŗ/�!��f�E]����,Ԑj�6l͕�8J���\2�J'{�ݺ�k��h]T��l�Z�lj]�ئ��ro)^M��,n���oo;p��:�K����
�*�$��XO���^�6n��͗#�3v�[m�Oli�B�G���j�B��WHZݮ��[�̦����.���*ə�������B�.ñ:�EL:Y�ub�;�YJl�1)�3w;$yk�0s�yZ�ۛ	�t�_e����c��=�*2Qכ�r"ѭC(M������CF��ۢ�V]�iu�(�j�*y:�2�3�i,���JA1dY�X;l���nt4�d��z�2�c��ǩ,D�a����Ѡ̥Qa}.��7p�ܥZ[��A����1��}�ug(Ǯ�f��+nΒ��V}-P�Xc�(�����!�v1O$[�R2�te���z�䦱b�Y�nn�w�\���&�G�%��ȫZ{�a���4\��G�D�:�tcJi5����ز���{J�<\�����V��sNg$n�]t�vrڅy���PL�0gY[�C���=��ٞ�>����dU�wQ���R=��:���t�;�YSk-S�oK��ю�e�$�d��*U̵��M\�fU�2�S��a�$����	y�͢ﻳ"Ǚ� �vemY����c���\����:��+{�5�;&�
Ը��x�"�d�rc�t;��M!ٵ�Y�ոu$N��H��r����V�S��4�M��Ӣ��Y���k�5tU�����oa�x;Hm��������ίD���dV��,�o1��[���vQ�U�2����ե<�f3yǭ㱛"*�	P���Yr^�ͷXX5"�}�rǕ�o���X�K��<��7igY8�ዝ�P*~�,ê���]��^����gy]EYL���8�/�0o��m��
��@���يsЗI�0�d�k@�]�k�e�Ō�+d"����9�7��(���w��v���&��F��y�&�.3�������]׌UӺ�O�\��u�mu-�wc[��!UG)]u��ۻ�Yu�=Ϥ���5�x�������o\�gw\��J4w�iK����9�ۡ���e��]v���#��]]��r⫽w�2���^S�����+ ƪ�S��+��s{9����W�c����z+����e=���N,K��J�ܺ�2����n����x�d��܄G��#��Y��dt�Kb��=���[YK�g��F���d�m�:�4pP�;$�k�QU+N��Vv9�/*�KySy�
�;.��d�� �{�M�n`��K��������@�͂=������.�<|��v���1\u!�E��7]�+^g[�]G,��3�&�Fj&'V���Z�b��u��& M���,f6l�.���aw�g�
9,���N�̉m��4�BB��Wy�ʻ�t�6�,B�+z�K֎��2�5/1���z/n�sl�����b�L|�E�|�'+�5ރ������Ss�����(��\���f��\��>�(�V�Sq�=�!}�Y��*���u{�n�Y��k��yC"�o�%�;�+H;��s�gsor��["�;0j.�^n+�՗cM��F������i=�++-�o��EF��q�T��Ïga���N�@9u�Zȶ�&ݼ�wمӘ������O�ُ;ct��y��][��,\[kqaݏ�@)��`�u׵3-]G�tx8��@Q�}��o�=k{}��-�S�b�I��-k��{	̦f2����V)�K�\�ݻ-��z�<��+��sn�ګ��'�*�f���to��Ͳ�w��^S�Wc mo,l���v��bu_X�%e�b=9�6��[��ޞ�LT�KFi�ԉ��xT�b���:��ˡr��ׇ��}�v&f6w%͂���.��.��]ػo���]�ge�뭏;��ud�h�œ8>��ٽ}�e'��ӣ8�¸�d���p_n���w@=�S.ik $�Ũv�5�֨���X�Ȝ�à���3Of��Wa{�70��sm	�3�=0Ap:��<f]r����K,{��{�Czn��먶�R�ýW�RVN��7���xnY�*!ĲH�]��:�X��u�G�Aԑ�]�y���\zO]_V���k:�3����ʕ{4�V�V휠-��c�n�9��7�*z��׺i1�1()���.��!XQQ�$�T��m�e��ؼ�(���ݴ�&;�F����ڷ����*]'n�l%���g޷�@)���I�k^���)�8����6ؓk.*�=۷K7J[S!�Nj8.�Ov�fVHz�w}�V�Ov�B����9�/o1�R������j̵�2�е�	lyo+��G�4�����5��ڈrV�b���+ka��moB7s�����`�t*���s k�ڛ�(:�{�,�0��R��g^vW`��c̾T��;v�h����b���*吃ocٌ�ڋ8�ʜ4��лݱw���j�zP�1�;�E"g�e��:�Y�')uA	��A���2�`N�>�ayٽ��Fƈ��dJ��<�ꂔ��\�>��s�	�����stUj��+c�����e���U���+,�~������v3
�v�}9�:^���O1��u8��WFzv��m��f���h]��v��a��Z�Z��{t�oq8/&�(�/<)��ìe*���idV����;�.{�����XԱٛp�f�ݙ�n��(*�YwDM�4�t���(V��$Y�pu[jn�Y���
�pO��oy>�O�q��,�u��;e�ɹ7�;ѷ�.�X�p�ʂF���P�n�l���R�+���GHo0�[7�)]ތ̹2���C�tգ3��Wdo��d��#���&Z���J���,�[|fiݗkF�r����ws1�y�z�h��DW֦.K:^�Γ��B����>I��L���i������[!���fCW��ً�GE���$�]V�n�2�غ���eAu�9(�Lٹ��f{��̲�3*Y��J\] X6�&��i���1a��\K�\bO�3c�7*���F䬩��z�]d���%h�^�Ւ�{v��h*�i�`�[�1����hp�\Y`�7	�)�8�#-��Re���w�f��x�N6�F��hIv��ۡ�̺�ò�+���l-�*�y�K��uoNd��m�a&M�����(F���,��J΂xʹ���j�7f�`�ݻPU�Ud�.�f�r�G.�F�I*��,��5�n<�ej��&^�ա���G�n@�d���y�U���ߎ��R��8i�{����<[:��y�����s;z��A綞 �O�wz-����.��巃CY[���mw{/��Aկ)PR�ǖ�$h�?F��9rl�Z.fwY2�t:e��}}�uf�R������nf����z�_��F�Əv٧�s�63v�A8�l�23�J�uwv
ܪX[��u�,Ͷ��"�s�lg`�/�og�����[�u��;�o��m�G�p�kC��������
�`XM9�D�QVڥ�e�V=.�������rƴU��JH�
�Z|qe�]�{�5��Ҷ�&�w������x��ӝ��q0��WO��J�#�&����;��J[!��*㧜Z��3�v�m(%��u��u�e�<��]������c���=����7�;�s:�Ri`n�[��ݲ���X���7�`���t��d��u���y\l��y2�K�p��(](�k�=��'�Q��t�K�=OR�v�[TU������vjr���0Rvt�zB��;�$��֪v�Y.��q�n�h���jvU�&�P�;��neңySJ��+z��#�\nQԕҾ���jc�Stt/���*�s4� 
j�4v�
إܑ�)Y�.eԼ(ul��)���q�z�)V�4��{[D�V��ݗ���]���V�c1R��Qۀ�h�٫y̩n�`�{�-�n�M=YȪř7p�O6��Y�̫tsLtJ��wy�;2��_
,�9�7����ORj^�90:�w�Q䭊묻�Q�l
����Zv�v�:N�j�}P�pn��s�n��&�Se���7nIG����w����qi��7+xfq�걦�CR�J$��Nn���FԲŜ<��N��S�
1R����-+��y����/��<1gx������=���'h���ՑBU��>].�-�����bTD�Ŕ�f�f����ؔ�m�6�t-}�6�y�&��p������<�e!s)��Ϋ��vf���`�hp|�T9x��oGs� �aA���b�6owyM��<n�z�a�r��{��� ��Aw3����Bm�{��,:U���#t72#u�ǘ���D���^�˃0��N��b�1gu�����怷��ه�n�8C�C���j�^uGN�2�)�]7v��U��E��&��c�Ԅc]����<J���ח��3[u&�RwS�Z7�jA ؕw6�N,�V:^��X��E��o���=t�,��ou��V���wwnaQ9&�r�$n�c�p�ב�bj.��F�f�,Vmm���ܩ�>I�ظi��l�[ �ˋd��`[�LB�.�+ojs�j�nq�������]Ǥ�N�G�h={4m0N3��W�N�}�{oU��8YH���$�<Q��mU��Y�����m�n��.�X
X������ͥ�n���YNu�;�M	���c���j;��,���C��k�k�X#9��������;�P*�k��Jo���rw��:Y�MZ�tr�w�iɧz�c��cq=�<�lY��ȕ8��U��!e�=�w�� ����@�1B�/�|�eǳU�z؛op�h�����	���P�<T�5�C$�휇u�qmf;.��ù{nՌ�wJ��[RB0S�yg�СwaU��Ywٗ��ݻ�-��V�v�V�堷Lgw������3�8l[��n����4��&^���V�^v\q�2���3�~�Č��95�J�'�Z��f�33�����/o���·*���b������cbR`��L��ޜU�z����S&�>]���[J��2�:�Լ����p<h��bmm�d+��3�Z�K���ɵ9e�z��6\j�2C
��ƥ뛬�Q�"�Iİ�9ARR�2���� ��x�z0`�p�r&Z�u��z�_]�ۚ�gm˝4ïj��j�`�ku��Ɨ�&evN̸���/oG�X����C����k��#�V믩�pU%�W�}�lM�hp{���o��&�ۭ¥���+�D���s�s;-���s��eXȐp^R�o�ޡZ��fG�ٛC�<���ֶ� �_V��'y��n�����	�7�j�Q�;���FS�هm׽F�tf>�\��j��tﲻ�Z�ыc���̺;�ź�����T�oV��O.��N횹:Ś��+�5nye�s�k0f���d�h���������:�U/n��a��y@�lf>�wth.kv��3�Ӡ��,�Dģs;���
e�Z�Uh�u��͆�`Vv/:�P��� ����ړ�T�k�8������X���ۅ�6..�+9�����Ǘ[�֗u�4��i���YvF^�{e�!�HҚ�a�_#%���neY�;Φִ�eefr]��*��=������D;]���]��$Wy�/b�����$+�ҷ�<�*-*r�ֲk�î�� ��k8��J+�Լ�h�k�V;t�_L֪�<��P>6�b� tl�ƺ��6��ޝ}%n���\����xa�v�U��/V��+���R�J�͵��F��3^��ɫCe�f�5e�s��j�/P[�c��rf�g8���;��A�9��h��v�69�����w[�Ӕ��v�t�"ɸ�~��V��b�*�L�=N��q�*�VZB�Y�W�tU�]t��F�K�<�e�B�*�Ŷ�Y}E��o�v:u���W1Y�j� +qf#�a˔����e��P-�V�g_�Tʚ9�:� V�<3��ų���L�䫩 �Q��ʬX��O+8�%3h-�#X���
7ٗ��X]| u��wX͔��e+V�5��Ovj��w�(�k�qAÎ]�*�SD�#y�E�).��O�6���ഋ7Æ��O�G�bYO�^u�x�;�PMh�xwO��懷��VV�ʸ�n8s����p����"a0�
��ps�t\��8e5s0l�կ�^�3nv�e�nSH�`=�`4���x���[��-�-շ[�Ԭs��l[����W�i
.-s]�=���޾Y��4�]C8
���Y}��L�Z�m��mL;�nt2c�;��T+x�4��]�Ǵ�r.�'�+���Hnپ����&Wue��ًr^��#�s{�Y�)�]
˜f���h�8iː7O+v�l�]�<o��%*2H�k���7�x^["�&:��-�97�%p��J4���kY]\#�sp��X��7���jr�,�JǠsuw���z�͂1y�;$�uf]s�b0����zȬ�6��QU��@�Z	}u�!��c*����ݕ��i�#���җY��cͭxj�<(�'�ƕ]1��z[Y�	�X�o���a�nެ�]�_e�׎]������Lx�8�>�ܱu���%��|�10bo�n۾'c�YN�V1����4�lr�ˣֶݺ�fp��tU��b�������M��R� �(���8�潀�t��[�׷�s�	V��:�Shm=��T+�\�l ����s9�qy�4�[sV��'2�;aif�ܱwR���@y*EQ,o�ځZ�B)+)JC��� �0�m.V'!bwgmˏ������U��\2t[�'y��}[H��]����o���h��7�v\�qV;ġ]��g[�sZ[�K�U�֥8���`���M͗˸֋�"{��u��["\,��y��!�a�����ؼ�m+uIg���w=0���L�5� 6N�ؽ��z������J� Ef��:�K�Veu�u;�T��Z�whŎΥ^iyF�a��W40H@
���i'�{X2ۖG�u̲ؒbx1WX��ؽ;O���U����;�<Q͠��Evt\\FT�Q��X��:��t���Ξn�R`i��[��6递�[�J}�#t�Qy��bȕ!gc���#u��M"�֝���Y��m�
�w$���4��[ǉ9�'a�d�.!�qf�m��Ky��Yq�ے�gu�8t��4rgk��œl�=�m�I]�v%Y����/.��aW[�Z;��*]KD���h�����%�6u��)���sxWLrf��+�X�.���Qy��d�ٹ��/�I�����+���V
{�Xb���N�)r��{��h�Qc�D��{'g=�Ι�/��
���Y�-Q�E��]����b�a��ѻX�N�q�+qu��%2%pqf�z�fz�Y�ƕ k�-|�E�������x�c�$VOhnJ+6�h���T��a��r�����˔�-�_!PU�:�E�\�X

!T6�Ju�p�.�-׏�]�ב�� �3�ٗ�h�o+$��L�r�u�yu��R���GNѤ�k��l[�OM����ٷ�ݽ�׃fS�I*�;˶�/y���Z�]#vtÕݡ	�1���2�]w4od���u���2��~����O���++���_�~m9_����n�m�*��s����X���l�=/�6�掶��k+"[�[�p<�Lq�suϳOV�׶�R�n{B����Ľ�ېD��.e��D���l�n��h��Ѷx�;5��N���i}k�۵I�u�{l��c��4	�Xa�l[v�r�^l�*z�[�vm�Fy�}[t��X9쮣��G�GP�O�7]�s�[pt�m�Uv�pc��6�ܗOO7+=����%�K��0�{�3NŜ�v��y�ˁU^���g��t�BWks�ވ8wV�}�n3�.�|������z�/LL6k�]ԯGAYy��n᭣�#�F�4�x�Oc�⪻�:;Nl�ƕ��j��Pn���0x0�X�n�6��h�Sq�sn-���n�=��7l�Ř���m��m۠�@��g�a��l��6��Zr��۷:��*��Ym�\kQ]O��K=�{wQ�N��NS���mõ��7�\���S�ı�q��n�o9���wk��\�����n)z�cʃe�ˬ[�@_�:��{fu��gG5�.9e�!�� �c�k��j�N���f1jn@K��=3ŷ\�Ÿ��7k:q�)���.̯9u��k�s�d�z�7WO92Ț������:�������:y�<j9��U�l빝��P���p�B�O�c��s��؜M��.�����n�<[n;'nD��f��a�g6�U/h`;3^�]ǻ=<9j�q��3��.�[u`JWG �������"d�+�Y+r�YPӒu���=�����6�z��]���v�c�^��㋬��>�`�lm{=ctBҫ�[��8D���%k�J
�=�sU����s]��ƺ��S�<�4��!�����k�۪��������g���p�N��>;j):-tuU�a�[��8��Ħn��[��=mn��6A���.�:�2�׷<��'��sW+������w�@�mϑ��s�k�։r�<��${W��WMb�<ˬ�&��&�W�/-�r�:�m���]n�� �;Oֈu���<����q{^�L�Xs���Ƌ�:r[O���0=��tv�1�z�k�:��Sʝc1ÞP�Ge^��GV�Qu�Os�a�k7'\�U�J�Wm5[.wY7L��s�Qȟ}z8�.y���kQo8�f# �������ɜXU��� 9K:IN;��	2�-]����a�g��[�:�¯*uԩ��x��FC����c��عN���t�o]��^���=�Ք@����.�Jl�-� ����GUyn�2�zϵP�Jj�ݽ�Y5�����e;u� �vJ=w��x��N1�V�uص�Wj����)�	�`�5Fnw
X�zf����lv�a:��Z`{F���#�j�Z�oE��\�� \�
뷁��'��8\ssqvj���N]ڶ�+��mր�n:2N���{�kۯg����4�w�m���� �N��[�6��������=�d��x�put�OZ��ō:��[/Vu�.�ч�;����ȶ�j��aU�st�����8��\�ȝ�ں��/<3m��%�q[�Y`��oNB�aFݼsع���܉f:��G<]Ng�u�Ыv.��.x�l�qM���r�e�c��j}��۫�ܦܑ�;]��Lj��oV��N����p�s8�F0�RU�綒�9��8�ɺ;tz��j:�ծ��xlH���j82mڸ^k�v¼<M����og��"��y�5��� ��rn8���˽=�`dۥ5�U�ۋ���uaz���� �X���N��^��`���]���m���7��ា.X*uv��P[rz񖗤�\8�n�����&����{���T��	�Z�x� �lC` ��g�x�)f�=�M����yݚݤ�ݺU܏;�:n}K�m�)�����u۲��th���)Ӻ�<Ҧޮ��ˢw[�@[��c�z�=�:;Wta�W9�j9��i!K�i�vu�mq`t�K=��9�c���p\�V㞸��lr��#V����lؠ4\(�:��ۣnjyG���K��r��^�:��t��Qu�;r<�^�@1�y�-�g7�^���$n�1��%��x�8�[)��x���F��B8�Q�7>Ĵ�a��
x�y��]֮��t�>r���9Q`���v�]v��p�۠��h�uι��w+V��!Փ���wT�m*f���\���q���m�oe��o��G݇��O]�������V�y�&2ք�����n�O]D�E��o;��]s�;]��u6��T���H1z����Lv=����=�m�3=�s�)�i�n:�n���kulsr��q�Q��ڭ#Z+�xn�\[���u��nl��@�����w<��-ۧX��yhd.G�k5����V]�ܕ���W���ĵ�8������[�������v0�9���n�LOk�Kj���yy����7����.�OW>[�ɠ^�D��� �'-G<�F��E�]��G�]�R#�0M3�Aq�.M�M�:�PF�K�|>:��;������q�;Fb�H�;	h�5'�¥+��s���[��dpG[tq��&/g��<D�:!.���cu\Y;N�	p�R�L���-���j��=I�7Z���ڋ��;g���X3���n�����M��\�����^���s@��1��`�83�K�z���P:�f��4Ÿɸ���j�F�5�Û�"��n���K+�����-�7�|���mOZ69:�Wnj�n���1О;��p�n���==kϵ�y�����\�Ì`nn10�.�V��[[%���a�ǚ�pSGd����^�uĞZ��3O��r�ck���tm\!�OGOG,����}@z�.�#����mj���z76����u9=v�hW��=r�:B��G	��7\q�=*�j;zV�ˁ���E�◧l��츃C����]^7�� �5��s^螂���WY0�kik63����[w5�f���d�S��������/Z�����%�'l�7��F��QU��a��8zx��G�N���hs�d'O����+��N)H[;b�Fn]Y�����G7vҽ��f��:H(ޮ��=�NKs��h��5��q��nA���p�{�����������d���Iǖ.�e䙎�3ɹ�sc{��;�\ά� �է�c֌qmf�X�s�I����U����=�p��\\��Ι�C��8�8v�=.��6����.�9��sl=�-�%�D�iݎh���/n9�l�sq6WiNx����'$�=��.8��a���M�=��m>Ŋ�%�1�踫]͉c;�}�2xx_]�Cq�cjA���g�<�%���K%��G3O[����mc�ٌ���\S�1^x�{l�G�=F��V�6��^t6�vu�3�X9k��A]+봸��F�9n-]nQx�C�w<��e.�>�j�s�y�A���)�)έ�tWU���`�E��Mn����5vm�����ﵧzF��:��)p+v�A{C	����mηZ�\뎮Q��`�;H^5�F�񕞷.���Ѵ�=���m��p�=��R��զ�h�JL�V�Ѭ-m;��;v��b�s�Z,ֻ�k�9[�̜�v��Gq���]Y�#ԡ��(hΠv�=̺�g��[�K�{�+�sץ���羊S��A5�/94���#�����Y���T�9l�A=��k;�]�v���r�ﭽ\TV�ѣQ��6d�ݺ�;��λɮ�獧3b��q�� O[�e��7qæz�&�v�8�!]���X��Z{5{���u䶞L%gvA��ϻ*[sF�e��ي\�E��v��U�'��:۵�͞թ}X�t�9Dw�C�w#\D�k������'p=��ݰqƀ^���n_K�����v�exW��7s�f��ǲ�����]�<M�6�oN{ u�����}�j9�H����Y�ǂ�t��M���.���<�mۺ�o:�mc&٪v�HCi#p���q�M'�68k�a���=2�v��6qh������upX���ۆ7:�#�s���ykx9NRN��o��p[��m�yHx��t�(s�Q��8+5cv9��|BC���ձ��ά���{q��;Q�3��<<�	��u���xݔ�:�u�� I-��[�`+��>ԝ�A����v�Ag�d �6lE�.9�1ْ�Q"vֻ[G/8�x��s��Vx��h�x'��=�'��M�!	���:nְ&����&�e��sG��n�)7n���9�x��y�6�N�ps��bN�WD�]]��ìON����ێ<tt�s�U������q�\�<�p�wq�k�I{v�u�9N����\��`��^�&��usvk�1��Q�@���]WO���8��I�X�6n��.�z�h���sA-Ʈ��1���r3�N�d#���\�4+�zm�^R�u�����T�T�W���Y,���X��f�ݻW�7c��s��q��vMg>��P���-.�oM�ۊ{%;��t�6���Y �a.Omۜ[d+�EN��x7�x��Հ8��x�7�r��i�ľ$e^X���\Q[�ss+�;]q;Z$���q�ܯ]/OU��bϻX�̓�,�-�����躁�88g��lp�pm��7f�u�jӎ�ݍ�5�+����V�=c��\b���ܐ	���q�.�]7Bn���n۱��<QǕ�����o@��޳֧��9���lFo=��ݶ�1M�s�A����g�[���uu���3���N�{lOk"k;���S�o,�֥R��஻n���	1��㧓3��6.d�uJ�r�4�v\[�q�[�b���dY�j�,uZ�0/&�7\�y9ӕ���v��ݛY�t˱�l]����c����!��lw^��Ŏ��5*v�r5�-VT]�X��d����D'�=�i6�K[���\ODvݹZR��=�U������ynlAtY��j�0�p��z���mȑ����g;������ܘ�b9���U�r	�b���[��n���l՛z��n�<^-�pV#��ҽ���2q��Okc�&��kIUr�N˲��܀$5�(�:�y�{u���rَ#�[#��t�L\���fD��q��y���cr�I9�qէ�v���@w ��;.Ū岩�0�s��Eԍ=�.�t��x�+Y�2p�g�u�c�r�]���d��s��8���Q#ڢ�e��@��,on�vs���u�D�!�<�]�3�nJ\�̶:�YB�V�rUܝ�w�4)�ٓn�s����7]?����������}|�w��hO���t�Q�J�W$��3�U7\���OA�X9e�^y5�-�j<k�lsGE��3d9 ��p���+��jKY��՝���쿧�pqx���+�A4�F�:��s��g�rq�Zy��S4v*�C�8*7���fE�q�m×��sJ��s\��낚��,�F��qv��,`:x���=�Ӄ��V�i��]�5��`%�lO\=we{��,ug��'ltc��ؠ���1�� �y��O������ؓ��}���ET~��>���_���{���z�Z�J�v����?��g�+�7���\�n��|�n)t�ևe�����G՗Q��®��fQٞ��?Q���[C��Q"���8�u�ʥ�;�kE��л����AG̧�GR���u���7�.�J�}�s2ά�K嵭9
_b��k��N��/��Yj��k5�6�5jͮe��U}G������(h�U���9%�p�U4�V�ؚ���:���¯�}��뎈�/3�lm�0���
�=uz�J�2(�L���ߵ���Q�X�β��k���ƾ�x�s3�#`�5��R���"�b�!����F,��k������n	m>���kB�F�^
cH^Tn�>�̖�-�!��2�˫&��X<�����(�����ǁ�6�yy��f_c��g]0�α�,t&mY��q��fBԄ6���+�V�_�D�&���[�<9�\�n-eL��4Gr�L�'V��u9�9�����t9�`S��%c��_�Ao��4�@D��F�C���(P`*���;��s�sQ��|���DX���1v#�cp݂���+�x �V��W�o,�;\h�+�����y�;%���2�u��]s�[���U�n��Z�@��|im�g_�����ʰ���PPF�>7D���0��AC0��)TU��]�o�?�Ţ]_7��@ kQ�jԪ\�4��Y(-�x#�[l*�$�ȒR� ^��(�^�����GZD��DeT�_�(B5P�4�SZ�XT�a٩�Ğ5���?NZ</�U�[��*�)
b#'LG*nσ�u�I߭���Sy�{1�*��yv�Q%�ܮ��g9��D���%
�\;%��"n�U���\�m����OX��k�Z�=�[k�����xɍ�fZz��
��٣e�%��Yv��[8�n�7���sс��:������l[�7S��<
���fOa{\])ث�S�ۣ&y�������ō��ۚx�z��}�,��m���-��{R��NQ�Ü��6w%��'�9ŭb-ڤ�nŻ�x��6��u�hk��umwly�0���t�N8��[�"=%�7'pq@�u�{�G��C��yN��	�E��Y맞�5b&�]ݶ��s���eպ�r�_gS�x���U��cn�������,p!�.�.�M��ݺ�ux�a����Ƌ���'�lnHq ��`���<�K����3�]����ۮ}�k��|{m��u��o�:.��un�c��r�6d�١�Ւ���[��ri�O��k7k�Z�3õp�@�<��n��G����8s;��v��tEs�YЇ���gK�����m�;f�S��=qHr��^��^,f���KWC�]�c<z�;U�F+���,���UK�7Z{����p8���h�5�W�p����F��#���hm�Y��7F���O`�����`ܝv2jhǷDz-���=p\�8���C<:g���\;��<F�{u��YZl�POfk��6�!�p��5��\�vz�:�����k�=�u7bv�SŶ�5�r�`��`{],�]���@4��4���#Q#����or!�ӫϧ�h�s�tXN6��oj�)i:;B�砭qE{O���v�Z�\� ��s�;�ul��B:��OG�h�^�wKCsН�Bʤ��[��뫳X��x�F�@Ձ����=��C��QƷa �U�)ź�듮�n�ͤ�l�C������՘�&ګn��hnѹ�[y1XM��'c���䳸Ɖۮ��2�v�L�tay㬖ᓙ<6��ǫ���pu�h�nM��f���5׬T�Ë�wnY�F����m�!���f�d��P��7j�}>�n���Z�u�)M�g�!�#�$�P�T�}I�s������*��=uh-�A�Rj�&��f��f����(	��h"���bj��k�D,r9�1hhƪ���0�띻���];��-\��p����/��Ӗ�ΖF��s�h�mGV�[]v\*�ܭ]]̖6�^%빨�ۭ�K��`�Pz���.4[�B`!��۫ۢ	BTQ�ƆN��ڕ��]y��S��n�՛y�0��� �k�s���[Z㮁���:�G.9�y�a�1���c�e)}����6�fi�p��1���.�ڼ�C���X�ɣ�3�n+�8��}�z�^�����E�PQnF����-q�U0��7�o U�%D�AP�I�S������y��=���������
A�$K��gNūyW-��]=��8֝{˭�֫PO Q,�:`����Ӎq״�sӶ�_総��|E�RT����~�ٶo[5��y��Ί�m��]Z�f�8:>%��Rd4�=��x�؎���o7���^��k^�z���5��7��{\��	�r�)<7
�.w=�G�[vp�sn.��^�ͧ�"l]�Q`��̓w�sֻ�A�mgu@�m���5���.�2�m4 �ƭ���^z|CUT�U1�E]Z�mQ�ESE���h�Np�%F��3G%��v�MSΪ��Ph�@n�U�j��$���f=|k�ް���[Z:�tRm�M'E�-��xs�1�{�9��}´�\��УD��,$�l7Lkٯ�>[{ӣճZ;�V�lg�M�/W&H&KiӧD�6��Yխv���wA�mn��^خcR;~VwZ���]����z�nۺ��t�W�fuZ�5�yvz��1%kCΑ�h:e1Z�{Թl��-���l��]b��Z��0�l"Qe�kV��)�N�;8�صo.[h��[}[\C&��h&�)2����ι�}��Vi�("i#�buY��J�&�����\�L5A͠�j�b")(��"�*��4�45Dk�{�]���߮x��巧�q�c�Ɲ[�ڦ����k���]c^��vu�G7������D"�ӠY�i$�=���ƭcv����`�\u�c=A�)�C^ �F�on�y:s�{[���8��B��N�jĆ��鍬�I,'H*eP~T�KLr���q�i�G�mw>:v���o��j�!��
l��M�{h�����{��K�V����ٺ:ĢA ��J�E��m��qط�*ӷ��Xݜ���U+�`�t�(�C�c���.��zx��Z�x�������Is&��j��QDli�`�kQEA�li��j�X���E��1QTW6��Dh�QRSE d�ژ��s�\�־����

���X-�[z�sӷ�r��our��_�8�
���%�ݹ6�zn:�g���e�6M�&i�Ź�����ۮgh*�6��v�P����[k7�׷��C�o�u�կ����k6�����I�B�mֽ������峟t5�f�)�N���&�H�t �٭�[k{�嶏o{N���=�޸/��l?0�u�`��\��{æ��k�ͮS��xF���
�Ц�+Ȧ�k�]c������[�`�����y�������%�J����".��"��I5AU�S�5%AK4��DUEQIQ!T�PDu�QƊ"Le�����p�y�qw�ڣ���6�mjq��v7������c��ͷ��4�׮�۳�W;ٵ��ۙ7Oc�Ӧ�a݂֨;q�&�q�����GX��X�>I;jy�h�s�]�n|�ۯ[F��
d;2�Ɲ��3˳�n����\�<As�+�X��S�����`u�_[�G�3R[�Q�7��=1���6cޡu�.L���d!�mY�خ�Xa��n��sg;	�@-ۚz�-P��9���c?R[��ݛ�Uv��sۭ��c9��m6�q��-�n����U���+)#���7{���L��q֎wW-���WM�aq�(R��%�i�	��=���:k�]kV���j�ֹpӶ��0�R��hP	5�^�=ͱ�9i�7�.:��\8��=�M�)P ��"[m3Zvi�8�ק�>:��Z�f��z�ֱH�B�S�|]$�e�[{��6�t�׬-�<va}��f����>�8��m�zA�����y�]޶��e�1ձ�:oV槰[���v�+c]d$H������x��9�ӷ��νk�׶7k��`E��	����O���G����B�B��h�*h���+�*壖*���y�DMEMP�y�I�DLG'�#��q�b&���Ӫ{=�ӯON|u��m��e�@�M����6��N|u�.��Xݜ��F����L&7D6Rc��{��=��-�c^��a��Z�!���l4���i�:�WX�z���zv��U���s��oOB�z�#O�6] �:[�X}m���g8�,t���mƀ4�̽����QTh�PD�t�C��I5�Z��u텼8iسk��5�-[o�p���)
i���ƻ���>|k��aw-;{�u���s=]�:I� [c�������߮;��9�ām�$�h��UEs��h֩j�USUSTS�bb�)�jbCY�
���-j����)
"k�3�ƨ 7f.����N0rث��)Ta$ߚ%�Z�c���ouN{6q}\8���pӯ{��4Z�M�h�=5���Z�|u���Ps���ձv�QRv���Sb�'n�u���K���$��wn
�u�+����F�Mɬ^ٴ�5�-;���`[]ǎ����k��Mr
d��L�I3\����v�����oK�u�fm	�\�)2A^ �Lr�;gV�z_s�K�|vs]\8�ΕԌl ���: �AMl״{���Ǻ�-k��ӷ�!DB��
Ӧ���ڛcT[*�pESSs��U�E�����������*�J��h�AEV�$��׏<�5�i �.�MӧJ�I5�����;���}�t�������S�@���]��O'MƳ�3n��3�����l:�-u�����PW]�i���;�����m���6�tُ_ٶ��;k7�綳z{{���M��d*!6�V�=ꃖ�/{�u���^�/��ٺ#M�TZj�e3�o�	ǎ��Ӟ�y��tֱo{b��L�D�HM�$&�=���V���k�=�usهz�Mxi�W$�4��
 ����':��Nzv�O;��3�'��$ �(��bj#Zf���P�4Z1UDD��U\�m���E�L@P�CTC5�����SM����������:�"�"�\�h�z�s�OU��(�< ��P�EΪ�����G��4qk]�������i����!��=�	���]�q5B�v�&k���;�y�On�v^8䛋�n�܆��lӭ��l,KV���{����N�x��!�],��؋�ܢ�s���X���s,�Hͪ��]YZ �̚�F��=����B�vs���w�u�|��y��x<�V�v%�k�Fl_?G�3��Zیۦ�����nj�n8����@5&C(���ݐ���`[�ձf�5�o�t�gr���֎�dh2�hQe7�f����֏q㷴�s㷜��Mxk@��N�TI���:��oC�l.��g>�-�6�k�x���a�4:�K�|v�8q�5�*�k���_w�B�A���i��5�.��Z�|u�ƹm�������	D�G@/"J��=c��^N����o����)���^l��3A��(�E&�N�TȦ�|��˞�ky��Gk�����q�uBO�yR�L�D�yk[���T)
�j�� ���s�����&��ђ�X������f�(���(�)��	�����*����R�h*��sïmoq���t���C��C�m��M����[���b�}\����o�N�={]�n2I4��B`������X͜y�G7�-��������RR��F�*M��:��\5l�ӟzw��ך���f�������+s93�u��ol�m0v��(�綁���]��}���G�7WX�M��~r��^w;=5�ރV���u�7�>)P.�)�@L��o6�fޗ��lӫ��w���UeSm�#E��ky�ٯi���_����`0:������F��R��A�6�+�/P�n�TD%�/�q����;+4^=ں�w]����HK=�q˙op�.�*K�9�v.�ng0��;��#,YR���i�;3#��
"k�s��d�%4��ha<{3b�^�ef�k���d6khˌ�i����]4�
�j�q:�ʙ0�<U� �n�ģ���mp���vb �Xec�Vk����uj^tE���Z-�6�e�i�ڬ�S���ݚtD��)�z+l�Q=�U��轨s{�TeC��u��v�x���^��Ry��v3s��dUꃘ�.��2�K[��e9IV2��~��YΣy��-К`����"�<�/���is屚�xek���x߄d��Oed4h'��[��]`�f��(��a��l����0�e��+-X[�^
��w,[gxT.�fRZ��"�@`�Pa�V� �ǘp�ڮ(b�����0�q�Eʅ�<�=� ��|}�rő@��$�@���&�5�r�FQ��!�&�V[~,�K���U��؛VB z�1O\��A
�[���ץcfP���׵5_Eՙ��$ފ^����gC�^ ��Q�����0#���tVYT���#�.P�Ρ-��;��WB��Wf��ڠA�nQ�c,�e!��7Pn;�Nq:=Ӂ7u�e�
Fr��n`ބp4*�)eF�(Bg�6-y#�IF�a�p�
G�r�u��6j��N�ݻ�����CL�6�h�ŝ6���1p�\��j��w9� ��b�!�9���4�TQ%P�\M���*� �=6����w;w��"��w��(��W�: ֤Q���m32�8�r��s�R^���+�u�.�,eh�9��3��s�w#��V3J�e�����oz�{ދHa�|�����ZW9ʪ��S4�x�d���w�Յ0]�UL�-u��K'J��;%�Y1�5Ŋ���#m��<Zܼ������q�¨[��cq;Oߓ��csn��x�|�	��4�{غUqq-:a�?��}Ӣ�x��{D�N���"X���H,:~ۿ�D��^0�RZ�X�ҥ���Hϱ�2�������/9�G)[	S����a��5YPC<V6M�b9ʮU2�E&��Xxw3_V
�x�f�m��;eq�ui���_v�gp����p�0�o��;��D�p8"�Z�cDST\à�(v0�LZ0T�6��(�b*���������&�8�IFٝD1Q|C�\I&o��>������G�g���ƌ���S)nz�LO���r��̨U�ӹ�Y�W��w�G�iU��;�����Z֝V�ۭ�������.� �T��Kf����������^���nݻP�v��v���5wE:/�v,*3J�8As���,�V��7�X|~��ʝ���XY+��xä�z�B�U�!��Ϛ�LC+�s�8�TXx���>��.s�0�wbm8m�[\�`�]�0��W��xy����r��D��P��[����3��{�prBD^W-	l�0�\�sT�ʲ���֙Z1��
���W:+��N�����smN�X�0��+]��]X*a�qqs{��LZWs��Z}ogiB��h� 1���O1Zh���1ERUD�476"`�b�)��b&�v�BD�ED�2��e�nCƊBD���w����ؠ*�U�����ؑ�;��1��[Mȼ�^"Ó���%s�Z�w�b�ں{�]]B���wFi�[���� :mĜ��`�6;=�����K<���E&ܝl�z3��wN8/^�@�J��U���y�u����u'�ۇ&���A9��j��]����}p]R�aI��g[��z[���	!�v��Ḻ�n����<sn-�qF���:�k��n6
N���{����gೂ}�8T쵋���:����7W����]Y=wmr�^�s�����^��ve]����>*�7�"�c]nz�L�e�:�\�*S<4���xoz�?7,j�J8��}XS�noǅs�\C+G'�)��q2�g��;��,9�q/x_�ڜ���Wc����X/.�;�.���B�ʪg���UA�W�{m3FV���6x8VJ�:ZS�(,9Ē��ΨU�ӭ�:�3J��JPE2�UU��wN��L�G��JGaaGjrSP��y=���2�UU���{�2��I�e"��-�����9\�;js��:L�[��z�4�;`�swo6m���Mq�A��9�֍i�nx�]%���̑vv��$��`��nv�0�V�T�ڂ)�;Nb�W8�`��qT0ex�6� 9B�ʥ��
`�f�g�tfzƪ��a���*��j&����TFƉj�lDL�#LU0��X481DATEQ�#�3ë��*�#瓾]*1$^���8�,K��ۑ��1Rؤ�;_Y�3ù/¨VD���T\�)��dr�L���Zr�*�b2��0��
J�m��C�qxVf�`����
PҙZ|�ꆔ��9H����4>�OUl���e�ua�
Eg�h��W��UcdަR)�%�8�På����Xt����tm�yU�667e;���l���U�6w2^�3<u\�l�n�v2��u[V�Y�Ս�[w�ҙHv��)�G�8��!�͙ԹŇ���o��H`�U6I�V!����xXt��u�E�%<+󚬦!�+-��L��^>N��+��a�U�4�H^;U�ޭ�>�1T,ei]Ϥ�>�8��;AUͪ�h��tQ�UIUi�q�QD��4�A�PQ-T���DPLPTcrO �G8*�J��{��TXx�7�N�a���4����|n�zŇL�_[��f��Dq{��#���*eC%��'wj��/
棺��뮧!`RGN����wgtPXx�WvoT+x���S,g�Ϛ��3�+�Y�Z�B�u��Y��c��m�]�l� ]KkO�9���e�;6nӀ��ՉD2 v�����a���:�P��H�j��R+��Z�*��R:ӗJ���S����u�V��S�.�xm9h)�U��v))����`��}�wN.(a��հ�,�;(����Ϊf��W��Lє��O	��r��|��+Fi��S0g��(�z��^>F8��(�\�:<�=;�E����>�0�󻳫H`>u��h�Z���������.Z�(��mUU4�QL���UADDMU5&��Ȋ"�����!�͡�9W9�~������zc�m�؄効��Hs5�_tPâJ�L�H�`�Tq{���R3�pLE3㋋3{�?�]N�%����-�Q8�ld��]��7i�;a�t��i���՟lI�{J��$�2Z���E��3_�VH���0eiߔ���b8�29��S��.�[UPtq�
�w���f��d���r��W����Pҙ�\�ެ0�w�..�.�����v[#dc��_p����ڻ����{��+
�8�:ٱYLC4����S+M��<�m�c�A��%]Ӣ�%�f��*�X�|�T�Lѕ�xOuCFr�Η�o�t]�y1��Yd�8��󩔆#��Vq�3J�q���T4�R%�
P�����*eX�*���e���墨b)����J�����D,A�1QD���ڠ��&*(!���ѩ���p�SEAD<l�RV+ybn4���ÇGd�n�s�gյ��s��J70]�62u3��9�k���բT:n;Ouf6�禧\�uӭ�<WU�0��ۗ��QV8�Q���k#��<������z�lGij$%o0!5�����sq6wc�W�w+5�����ۃ��z�v9��cZtO�v�Q1����$�0One�S�pL����n�bۇS��]���l�|����㫞ߏ{���}��,"�`�����uQ�����9a�.o8��w��o�4�Ω��^������(��l:����4��*,���^$��(U��>u�UWZ1=�h)�3�D�U(:w3��J�-����x�sgt�8���x��U
��w#�UZWs�PP�Ua��W�y��ET�j�WtTXt�ԥ
��#͊���s��W�W`���|~�w��<,:;�m�B��Ay��c+��I�-T,e"��pLC+�q��P�)�\�o{
C4w7�k����7`����0�wvw)��r���Z�)���U
��v����/��������tU�DI+7/8w��\Pãl��BwPq���+n�7h��A�%�UZUd��;��G3f(U��g�N�R�d�Õ�C>w�����m^f��Q�J�V��7n�:�k�i���b��K�X���s�(-��QQ%̺*�b6��UATT�1kA4[D�*"j"y��)��x�sǯ~�2�V���Z�Z}ogiB���3O�i�QO�8��������W~���'���UU2��ʹ�S<>�ں�T��&l�F�#�!�A�m���q$�'s5��L�n�訰�$��
���*�;V�QL��T�Yњ�r�[e-�K)� �_�ߧt�LG9�d�z��<G���e"��7�æ�s�_����	�ӓ�N�AG$��8��h�x�X�t�ַCy�{f۫��ی���yi�-�� `:�}�Aa��5|(VG[��Ҡ�iMI������񓻷�Aa�7�w�㳎J�%T+Fx����L��+Fiƈ��X����oV
å˛;�\�:�FkVFث䄧m��0�ݫ�A`�ﵮ��v6�p�9�bÇ)�j&��)幵�s���RS�@D�Q34SMUQQDADT�0�	@�RK�d��Z.�xy��դ0]�u(�ѺA��$��`�Us�;{pP�S4u3f(U�G�'|�S4g9U�T���YL�2ϩ��Uah���_p��w3Z��S
�����*����<R��u�-B�XxK��fj���9cl�����x,��Q��gt�t�
Χw�qۖ�0ls��
Hev�X5d����a�'fog4�4��8R����ӛ���UPE3�q|��]0���Q�h����D�ua�+Jr/b�W+�e#�N�2��i&l�P���{�UUR�g>����DYy ��U� �^��H,:~�p�P�9UUL�٪Z�h��X�v
�|~Y�笍�9h�+v��,9ʪ�d�z�X3�_S��3iX����<���1�T���� �#�`"��&���0E;
��)))� ����&��*����A<^�������$�5X�ܶޭ��&*���9�s�Ԙ�c+H� �VS4n+�Z1��S�;�������o)�;L�N��̝c�����qVXv펣��מ]j���u�S��x��V���c<W�/Zf��3�SL�_y�q-L>6f�.�)���rk+i�c�r�V��0^w6wD������I�c4omN���<W�'�P�s�^0�L�y��~��V�nW� ��.l�U�D�<*fU�S)�M��Lş�y�)�>3)�W#*����#-}�tÜ\��y�{�,)�����CsN�6Rb)���qf˥P��4�|�U�brU#n��z���~N�ꆌ���s�֡ZS�juB�����61iL>�B�U��k]k�,�����eX��{�����.�[�2�V�q=J;"M����8�Z2��  	B�<�t�W�u�аn�G�2��q�x̀�4­Q�!��N�1R��[���-�N^���EX@H���3"��9�sO-h��7M^
hb�13J�v�
y~Vn	��FX�AB��q*;MO�\J��}(�f��o|�%���t�b��KPx��v,(yo%-��X[+㣗���iS;�����G9���@?�����X�k��I.�a<�V�2�i�Yvf�2�j��6�DU�r�B�8�Ӿ�P�ܜ��*O��f��̩�t $�U�ؓӒ� %5����丩�-sy�Y�Sv�]�x�ޔ��1�p42�ʳ�V�+�-�+�E�x�:Oh�i�~(gcJV�:�7X%�T���R�W��j��pVin9�zQ���-�
����Rhkt(f�X�T���*�Gۦ�6��z�Qv�[!�y{;o�:(�&�����=9�z�X�����/��4}�\�E�'v��3�^y}�C��缥٤Y�F퍚6�CCF��S�  _#ի��I*K/=ܧG����Pƺ���r�4�y��^�H��SJ.�V����7w-B���Q����ۀA�CB��>����~Db�!L���I��D�S,��)�����=t:��F��B)${�sMP���cQ7[,S�oͲ"�J���Gc�l�oz��qXV�m�XI���z;d���3�\Tjƒ�o9�Ƨ��I.}���ȴ{<Z�7cq�6�'g&V����Uۣܻ%J짵�qk�ϣ�����
��l�x��z���[աG���[`zu�x���ד���c-���u���tG/��Ϭ�Y��w/��O~�}��i�9غ眯mӲ���=�-V�X����j��ǞA'!A�<W\��]j��C�a<�ɒ6i1��^[�y��M�qt�ܕZ^N3.�D��(<��ڸj�&�����'�����������V��;�[�ɵ7]y-"K�x���PZ٩�6ۗ��Ǉ��P���M�OW]�Ƕ����cW8����\rc���5.����ѐ�O\Y"�]uٶ���g��L=v��z�7�rl7N*�;\�F�6��m���cW�n$�,TV��NH��,s5/�96��u��B�����G3u/����ql����5t�kBn��eY�������{n�W�Dۨ2�ժt���M�i��3Y<�kOܛOg����I��V1]���y�ލ�37U���� /7Mc�E�D�kr;v��`�ុlF��ۛtK]2���G>DD��\����2/7ƣ��y�s��Y��MW�[���tt�����n$�;����;82Wfl�/]nn>y7�J^TT胓����x��t3�>t#��vnm�]tu���ݘ������d����ץ�Bi��7f��w�\㦨皇96v�\����	Q�Ƭ���k�R�#�n*xs�;��mb{mz���7[\u�_8��a��SѢ�fZ���[f�����}>�-�h��suj��b�!r��:v
� Ne�
vu�^w'��6&5�� ]7��=:�[��`�1˲s���1$q�ժ��ٵ��8�{4���J=�GY�^��{�;�q�u��:�q��d��͵�i���']|(E��혝���ŵ�f�v.��Ӿ��j�s����z�g��Q,�<��\��xU�{ �����ȹ�B���8˸8䮜��ѓ��:	�}����Wn�v���9���;�upOU9L������������_~��5hqTIMPR�V-!��r8�DIr�D�4QDEUDQP1TTՂ��PQQSۅ�T�w#�,kLj5ɞ��4s�ټ�P����8��Os�%�ۏ�W.����Ż<�Ǆ����)�����d��g��ә ��q�6*�]�k�u��KI�ǭ���.�<c���{�z�v��;$�X�^�ny��ɳj�E�m�||u���3v�c=�����f�u��R�]�^�4�W�v��>��OT��z"Fwͻu�x��S�ф�ݱm�z�:�T�Jv[G����^�;���i�Ɠ��e�ax/-��6r�k�Y���k���k��9
��G�/C�Z;+&������¼~Y7��Lӱ9J�V1���'�*�.s�CE�n�/t��y頛*%�ʪ�9Z������<a���fEG���q�8&r���S>6j�6KU
�Ki+��S�I�L���r�P¹�WZw�%&WE��ӻ��/xK;C�����Zt�ŋ�T0g9�W4��8R����>u7��x�ruS*�s��s÷�A�{����R�T�v����s7�&R)�9U�s�>�2�f�ϝEҡ�M���9�s��?w��DU3O[��`L
rKkq4>�5�/'��k�=Q�����AV�]�Z6�JwH,D9c4k;'U2�W���)r��sJ`�l���
s�;�j���U�����wL<S��O�#��1$DD����T4�r]�mq��(�H���j��)�H���*"�h��SLDX58����������W�o�_S+ĵ!JS֜�L�8�T���b�[���I	iդ0Ӎd��c+�y<R�"��ULCFI;���o~��0�Z�F��++�I_p�8��x����X|\��J�X3�c��T0g*�ʤV|�����ɬ^�ʤ�6I\��ਰ�R�+i\�9��[�e3iR�P��tŷ�{�9�q%�}���).�GQ��n�\��ۋs9�γ�"�y�J�[s˴����:�v����k�S+F"<�1�V_�	�2�cs�.r���H�x��gi2��:��]�+!h���o`����Wt�J���V���P�����B�g�k�_V�.s��xY۳YH��J�tR�]�(X��)�8�<����\ERDD�lj�DQL�TQM6Ƙ�cX���b��`��"a�	��1DМDCZ��y���h��^n�wb�X/���|�9DXڮ�8�e2���^�1S+h�l�P����ꖡ�(�s�ω�2ҙ����@
��(6�}�/���J|"���7�֡�2����f�ίw�E��\�9W�5�K*�����1�9��`����j��٭���wh]�k#�r�(7��Em��J�e#��XC�f˥2�v�b�"��d��ʮs����]݀����<j�Hz��+X^��pP��^�u��s��S^�R}D抙�+JϜަW9��^3���;^Q��n�Z������{b��i؜��,�*��E7�1CJei���� ���=���Z�t���V2��Uh�c��2�S��1B�WO�w�/��p?6�)���FvpEm�!�"m�UF�;:"(��"��ն�
��*�E;ۯ=�wo����q�eKa#�^���⻎N҅��ҫ�\i�oTL���JT���u͖�2��Ur�����(��s�ε�u�]tJ�h��h������]j���D�h����s��%ۆ2�Pѕ�QP�)�6E�L����a��r�c<W�4�W��/��k�W-��l����.f�Xq.r����¦!�������Zr��\PXt�߆��QQ�P�]eX��Ih�X���.�4�UW�اTL��͔���)ö]eA\��۵�a�s�.���p�õ.	�e3G'�E
C9ʪ�$�ۮ��x_���Ū�F�\p�ڻ����P��*����`�KR�Մ0])���!��L�&q��\�QTD�V�"�����l���LD���TQAU� ���������z1����	��}v�2���tc��^�+��K\p:8��7u=k������T�-��l+bz�:��0i�Ӡ��<۾��Lf9��t��k���/1�k��u����ƻ0�]�Ϯu^�_*���=I�$M�#%�;�30��@(��n\�q/rSh���v��!�[��ln�Ku��q����4j��m�Q�snX{p�Ov��n�8���%���Έ��w��w����-�t\�U�p�t3���q��S�4�9��`�"�
�	Y{1�0^�t�ݛc��N��f��*�_��c4��YLC<Wr9��UUB�eh���CJg��T��J7cR��d��`�a��sgV������|�JPѕ�s)B��xo%�Z.qs�?m�/�S�%M��΅A�R��2����LӜ�8�5;7���>��J��+Jnw�Qܲ��N��+���s�������C�t{�)B�b;����P���W4��D4���]o�GA��a��xX|l͖��c�W+��LC+J�|ࡆ�˛tTX|s��f{l"*e��^碲IY����XC[��{G6������m�k�`�4c���[�<�ޯ\�g���3�Z}��3iMd��e2�v)�$��Xtܾ�wNtæ���=\r�N����Շ�����]�����MEP�O-r5UQTAO,�6�CDKEC@��PL�ptEj�����E!�_Z��)��払�<`���K�7��J���ʑI_p�2��l���3�7�G9\�x�I�V0_;wop��tߏ&Ԋ�n;*�n��Ĺ�������/b�4b*<�L�W)5)3
g���صC�0��5FZ�Ղ��wz�U2�W�W+�OwD�2�v���8������>9�qj��m��%\�HxH�J��^:��:w�,�u��H\pU�񋹛P�X�k�샃ꅒ*;��:,:3J�$)B�sO�E�LҘ���us���:n�l��.���S�;��Z}2��yi�exnw��
�sJf�=�eh���J��u͖�U�YL�|״="�6ڲ�"�gt�ã��_t�0��w��V�9�
6�+P \�DN�*��"i
9�TAT15�1SAM�P�6�#�qq�¿��;�L����<s��u�k,���W�IN੅W*�V96��<Ws�8��9�q�
Xq.x{��բ�2k�����VpnJui�����S�.$󻲔*�f��=j��d�.C#��=��~���	��"r�_�evǓ�z޵V�-Q%��<��9zՌԅ섇v��W��p�u����w��� ����R�R��+��ʪ�h�ұ��I�b���ߠ�rE�j��gp��a��P��,b$Փ;�X�*,����7�N��Aa�+��UV��d�t�f*eh�g�oUA����&i\�HjK�2��x�|�	��4��{�FТ�r��N��.qtO;�;����$S�S<I��Tʱ�_U7|��WA͹�0�6��5��&��cF�3�`������*���X����J��g�E����x[άꂉ�%��4).be��|����㜮g���Hg������c�.�0g<W*��J��@��c��tvN:^<�	�0i�:\W���Ϋl�rn9nc ui���\����o8�e1oe�e!�}se*���W֜UT4ei����
ҙ�s��|����Y��:~�w��h��R��T0�R"jRf�1�I��*a��m��X��E�S�O/��oS4ex��LÜ�b29��a��wsWy�0�n���88���fgT,�UW<7��4�#������5:��g*�ⱹ���W����"m��A�9+]�tX|l�軂���r�͝AL���jLL��Zdk���un����dŬIl��Z4PElhJ
��". �� @�!Ƞ���qM�]4u���s� ��dxwV@żyQ�;G��Xݷ��r��8�[i���)�A����<��n`�%�;�:����	>��j��nSW2(��Ƴ!Y�r�񉧗�\���﫶̌u�Oc>�����Z��4뮄�c>�۞C�vlf+f�����/��lq���G>�A޺�֞�=�~���vZY��CŷG�y}��÷<ga,��=4��҇���n�ǻ�׏��!�M�W^�;����Z�� 9r��u��;�s�u�r��cp�tg��YD�x�X��:i�w���ZC�WY%�X��.l��B��"L������Ȍ�E"�4�B5$�W8`��;�B���qϝAC
f�oe��#��ޭ8���~��٪8W[%w�^w30ei�)B�L�R�2�\�g��N�t�h�Tq{��R2�e4�#�mvH�R���E�\_����B�b;�8R�`�ҥ�^0g+�Gs���S�x�=���mI
�N�IN�V3F,�P��9�u��(X�i�
uB�g���*eh�Uϩc���.�n(M.Ϙ<��ϖ��7n\�V�u�ղEt=�v�.T�����9�ZЦSWx*f�V[���2�c�.�+
g�jB�+�
�����4����CK-�n�l�Igt�^2wv�N���5�Z1Q�Ͷ"kZ�w9�Z�Ȩ*��`��&` H�N�s�T��٧V�x�����<a㘦�otI(`�<�QD8��7c�v��wE�a�s{���)�Δ�r���X���W��^��,>3�ro+"�QYj��t�s��IJ��iϞl�Zc�.�+
b�_��otPæ�|	����e�H[�,<a���wJ,��J����L�z��<e�PT�^9�W���7�(Bq���n	�8�N+TKZ���(����;aql��+���+��9wR�.�[�4�+�0^w6wJsnj�*�x��s:W9�`�-HR���Fgvy��%�ELr��p��ٻ��2���&OZ�`�Eg����W����%�,>,�m�AD�B:�:�X3Go��3J���T4�QR�ߒsR���{j���zsߪy"4�%�fP�7\n��e��o^8�-���軮��V[Yu������t;�x�����>��qq:�7�Y�MRƻ&v�J�6����n�P9��6*1��F�J�)i�ù���j`w�W��:��e ���pGM7��܄�\w�`�z凗Io��>I��˩|j�t�"�f��'D� �[٨�E�^�#�f�����+4a��K������[�z�S;k���Ud��2�im���挹
�xI��w]�o�^ѹ[o\ۥ\*�	���q<���cj���_�K���P]��f���c[�zL��r{D���Y���=ȫ<dޔ��4&���C]��W�f۸Eӌ�����4N��t|�a�7�\5�rv&��\3��)�d��XΛ&���J{(�#<(����ڑ>7R�(�yL� 4��2(]K(�rF$��E!�]ݡ��!�}��c�P?hTՏM(�����bb6H|�t�C���|})R7�q�f���� ۻw����/<]"V��ʔ��DpWn�.�,ٸ��oY#)M�ˤ�ۦ5!+:��c��0��M�CRc�n�Y("WY�2�!ڧ��X���V���E�ܤFV
w@4�.!�EA1Jƅ�k`�kn��,�7�w��ѣ`:Jԡ�J5*��E_^1ӷn�A�)a�8�t��]h�3���/�[��͝����X�՛��`u��\)��T��w-e`��D0����Mֺ�P����>��j����ڵ�ֹ&�M�LE3ɭU%DQ4AcW;���Uy�r�Lw��(YLG��V���7�B�cnF��}ZXʮsJ�'�J2��E)2�L�9�L�2���qyaLш��(Q����n@nW�:aχ����8�NZ�VӿM��b9܎R���8��ݓJ�)U�7J*����M�Pj��:����[�nD풧��,3�yJ��<z�5[��"���iN訰�}�wE�'�aPњV_���aL�mΨQa��wvH��yBGUqӫEL<e�'3��0ex���uCFW�3f((,:=�j��Pâ�߸��	YUv�Y|��Ҿ��
S+GS6b����#�s�T�ш�抡�+�}bv�l��X�����:`���su��
g����e!�w"�P��W�w��U5Q%Ru&�*"��H�jJ����������A4�����N�xÞ��H�Lh�̮�yi��!�s)T+x�r��pUZW��D�^2d�e�g�r���Bm�,
劒��V	����+�q<urE�\�/m��95�[1��q�����Pu��%}�t�⟷}X����7;I�S+Isgir�)��|੕�3=��#%n�[erӫH`�/�l�
��ZKR��VSٓ֙Za�����q%L:/�o�A�Z�����n�,g<c�-2�g���B�\�g��=�T�H���ѳ$G�H�'*�[N�,9�z�
C4�չޔ��w��)��4�4ӺAa����j"�YHdr��)G�/Z�h�Er��pL������3~tTä�D ��1�N�*�(��F�KgDMQATαDEP^<ݎl~��-slS�֭����s�]��뭬n=H<�����_o���(��tn��<E�������\u�l6��vp1�=F�sϮ�;*��r�'M�:�u��=���c�}�x���G�n=��;�&�Ŗw�T�p3��k-�1VE�:;kq�%3]�Q�D�� �םNsH��'7m�鴷��u\:����9�ƶ�%�N������lמu��p/]��[�EOcu�'~��������p0]�{y�Ǉ�k���iͺ����|��3��n�wmn�"ЛQ�d�8���?���?q�ws���)B�ei؜�)��)�U\�,g���`�'�ż��§#�w�fZ���c�-3��)�"�uB�f��͐XS	��k�.r��u]�Rȉln�*�JZ��E����X(`��h�W)�8�I��2�K�;J�O�}р4)��%h��ࡇ+����J��EG���e#�{:��Ü^.f�ӝ0�����T�aP6�e��Ҧ`��RlۥZW9-H&U��u�-2�f�<��¡�4�*&�y�a���ֺ�r6Na�on+��=�>�%���s:��zꄒ��A� !�K�v��3�y�)���_��)��ruT*�x�/Z�re"��7��exoz�����c#]�S�.�����p��y.�61�b�f�9�U1QK\؂���'�b��!��^����߽{����������ukcvJ��Yb�R��Nb�`�ұ�R�,�S+Ĺ���e1�S���x���A���jG{�o{E�L�'�~nm�����ަi�{ܯ���H�?�*�0���u�F�L�۶�J`�e�s��3�q�/Z�h�7����4b+��)��R%��w�en��۩��]O�ۚol�;S���N��WG]��nw!U�0�c�{k�����L�N�3�3N���T0e"����i����gtPXt�b�[QV��e�xVnoA`�0�_�sE�4�W��E�PҘ��IJ�\ў%I�����9k�Ӧ�w3_p�ù��t�����hm1}$�
H�X�����j����M14PQͦ&���7�ׯ^����&�q�g�w'n�^t����\񓹷�Qa�!�تc�c��3����ꅌ�7S�1�v��#�S�(,:_پ}Ґ�����])�3�G){�g���w����`W
�*�z����2ip���^��/!��;�������$F����lv��XW,��t����j�c4�y�4ei֧`��U��?m߅��:<�h�9�+$���9�
f�RE�L�"�Hϱ�1�Iz(sx�s�3��R*<%w�T�Vܖ^wJ`�<�l��I�*�U1=��¡�<SY&Re���ά�q7��جD�RY�<,];&Ψr�"[�C#��S��g��J�������0�:q	UA���ܱRWJr�zf�߅E�����쮠��nRv�
C<w糴��3J�w#��e2���JPE3N��P��*�s���к����;X��f�O/!spF��c�u��hz6�����+�Xӣ�޹��.�s-T4ex��;Z|��P�)�#��U�R���)�g���_j�%M�գ���<,������KNR�U�GrH*e��+.9J�0_�o�b���K"v�tTX||�'�B�b>NoirUS<W�6Zf���͝ҋ��G�F�xR1H�32�B�er��'tU^+&�1��8&R)��Ϥ�
��W\!`��L�"*�[z��釅�w�5�<3�s����&aLG�'�T+F"L�j���p�[��B� P�C�U�4m���hi)6�U	�i�b�k���`幮�b�oF��V����{e��j�6�����$]���lޭ�sۣ��.�񺳒^3D릲������v�]lUw>����٨���������WBd��@xLUZm���ィtq���-��6dm&:Ea��tm�n �v�b;�����m���z.(:.�\�j�h&y�7fNy�`j���-�;Y����x�A��w\�Ɠ�HxG�t�z�5���^��gwדp�뵷3��tŐ�ة�S���e�.c�-v����<��7��P�H�UU�[-}Ӧ���8�XS<w�)�[�H9U�ɾ�� �]?g���o�U�M7lPE3Gi̥P�V���UZS�/�|�z�9�ӌF9�[y��˾���u�Y���!�)ȼ�PCY8Rf�9�M�t��3Ioe&s#?\Hkcay@i��oVÜ^N��Zw糴�H�h٪Z�h�x���ݢ�������[]��Z;_Y�2��M�f��X�R�V�z�2�SN^��ex��zu�U�ۆ�ݶ�W^������q�<���
x�쵸����=����v'���Tݢ�/)2��i֤�
��tϜΕ�5�e*�������("��<;R�6�	]p|,�V��ߧV�9LL[�ʮV�SN�A˕QC%EM�5O@V����b^1�oS)����eWL:<�hϹ�vK��ZS���)��9I�s�D�*
��?m߅Շ�E�����U�Zm�e��2��l��8�e�:�X3�g�j���W����&"�^>�]!2̑;,hvҵk���]Z*a�UKs¨`�qړ,ei.l�(U�Ή/�x���pq4�ZuW-���Z�[��ՖՅ[��P��;v^r����/A���c��F�v��a�2���0�J�6Z���F}�
��S<e�;J�Xa���'h�UW%�eV��xN�%�UX���s0�4�I��h��۪s��������kln��F��)��y/��}"�UB��>�ǡ[(��"���(��E�$@���|�.v���;/K�ӎ��;�0^3���kj�:���ق�aL�V�Ԩ(U�G~N��LC4��IJS9�;��e1�ok;�N"�TA��wNtç�غ��W��ިh�����LӌDQN�U���[�E+��rG	K�[Ïu�^"j^��,�j�y����m�7Bkmzd��d�L%��^�,)���n�� �^;��P�br�9
���IP��9�,o�i�[Qd�	m�Ӧ�v��B�
g�3�:�V1�qYL������]7��(Ɯ��`���0�h��ުe!��2�2��2�S��)B�R:��PG��w�����
�j)�0K�)7t��|/�6qCFq>���S;�t}¨94�Pj�A���Z*&p8������}��E:b��EP��nG)ՇLD�f��L�V_�qC3�RoiB�f����3F|q-](��7F7�:��"*n��=Rs�a�rѺ莤���������Mn�O0Ғ�!,M�"	m����j�$�.�B�f��I���3Ncb�PF�a������d�ZQ�otTXxϚ�P�C<a8g!�<V9;��������s����`F���Q��Gw���c�I��c4�rH(YT��uC3�y/h�JMW{D���uGk#D���Ë��3~}���m��)���U
��猹!J�c>9��G<�NX9b��YJwJ`�;�JLÌҹܒ
c4k-�|��O����X�c}�T�Y��ԩ���W��|.�Ge�ŎL��E,���b:�U��HI-�o�^����G�7-V��&��3�����u�kAΒs:�
����d�>r���ڽ{ �]e��*_at%;���\C4PS*%�������

�kF�MQ�P�>&�v��O:���j��%ޢ���	u�^���g%iY��b罱�8h�l^��L.68;8P`����c��7��q�r3C �E���'�Yn�(�`#Cn�P��Y�+Z�o ��o^�q���ډi�م��x��y޵����mWn���5�o���fYm&��3d�+G��sh�X7��F��:j�]K7�$�QW͎2ژ��
�l�O�+��qQ�F�޸h��%������|uS؍46"����ϥ�۬�x�Q��ɩ� d���ԫ(h�����v�2��]�OG�^Z���h&z�\S�0�'B*O�Ў���%jܬə�!�+u���խ��^$���R���jW� 8�o�*�=r��b�"b�#��w)I���a@[�kut���.�4�t�)Q.PLG��<�$��Zt*f !5F �X�R'h{x3,��*�(�9�C���p�ӥ��kGX�Q�sGL��b�z���)%Y�9a�9o[]��P���3"f
���{�MV�DR�	����e;7��<膸Y�0Hmܚ�.ǅ��5Ab�(ƦC`f"a��+"����:���W��		\[������c=�h�5w[ۇ�]n�on��;v�g��nAKA�]=��YZ��vYpl@��=z�ō��l��Y!��"v..z�7!i�qf� Rذ�!�w����#��4\=S���0VY��
�nv)�em[�:�n�F��նNKsq�W�Ҿ���p���ی�J�V%�yz�i �(f)uFg�U�"��JrZƃ��w��l������ r�㵡Ǵ���tu��Cԕu���F�n��son��:�M��7[��un"���n"X��ɧ/9���s]g��9�4�m���vaV7M�6��7q�n�c�\�ܕa=�ngCj�;9��.���rb��]�o9���rHۖwh�ŧ����t��=3�F��X���9w8۝�˸���w����i��7tΝ��&�EG���2���\�d�;#�sH��t�ۊux�>�*yU���&.E���q>`.t��^c/������\+Ż"ϱ]��ka{q�Z�Q��.Dݱ=�آ���^2�y�q�m��[��Z����d�<�9G �Yۮ^�}j�1�h;0�g-crqƻ=����Ƃ�9�\��[�9��y�n8O,hگ7����ҽnІ+�]��t���v�us�<�i8�ňnuН�q�g�^�8��\6;<Gnt\�$"<����pTQ��$훳<\�M�n۞:��g�A�;v�W���q��x|�ĶC���ު3�Ҏ�Z�9N���<�n�]jul�\mc��^�pn�79�3�@���;I�t��@��rI��q{t�lr������z6�/>�Ln4l�ͽ^K2�Ǫ;g��tr-7:��5��ݸr�<ݗ�j�*pC�u�j�ד�Jq�L�Ft�M��qC���6wZ�U��]���@�ȍ�Pf�"m׹�>�rQ{>FƦC��Z:㱻Nn|K�׷O��m]h�4��N�Z�ouaݷ܁�M�8z�
�́�����m;���=<:�N�
/b:Ʈy�B]h|���֞��2b=1��ۥ���FTЩ\��g&�q�����O�:@���Q��wQz;'X3�v��=j�j�*���n۵�e�#X==5�\(���Pӣ3�T�lQ1̘�l	m� �GG�����m��ŭ5ӓu7�q��{eܞN��l9�e�y/h �y�s�Ä��%m\z���V��]QXxx^z��.8�`�[v �F�5t&��}s<�+�`��G[*v㮻Fz��=��\�fw�⋚:�9�ص8]�g�n����:��;7:��f��8�8�=��K�[Vz�mP�����B��=z���=8��՝�\��:�b��]�v�Ӓ�UÝ�߷�?|��+�Me����8����ӹ�*�)��풅��j��z�r�ݖ �c�i'F�&�Ѕ`�w��>C�.��`�Eg�oUS���蘎3��ST���	UN;���S3�N�Hf��l��vM�P����D:�Ix���.�m�����t|n�ե�����Pѕ�(�S*ʦi��;������L>���D���IE� ��^��N�E����C4��Ϊ����+.9J2�c��ؤ�;Kku8����å�sgp���]*1���Lќ���{�E����Q<F�ȡ-��T�A��sޛ`�i��wmf�]�y��5����ݨ�{D!%�AYl)H�t�0�f��K^+>s{Jex��R�31Ә�T���R5����v7��sHa�<���T�n��+��$�5�4��EGU�'d�
��US+�:�֡�1L�9�^�W�r*p��FQ�3,��]�S�F[s��XS<w糴�H�4�O�T4f�ߔ���sIp�e����$T������L�y��r�|~�.�T4g�49���s�>QJL�)�2飲
��i�[Nੇ�f�8���l�f�6wE)�u�l�野/�7�����Ym*u����:g1���8�]�ԩ���1��ݻX��[�xj�1�����z�������X��.l�(Y�!�S)s�������i:/��Qz�VKD�U�l�3��nu3��3�<r�C�3Ó۔��0��Y���	x�|<�ٮ}P��;������1�'T*�hܿj�Co��5:��Ab1E���W"�����Mp�v�U���+�A��Ƨ��`�ʉ�$��U+��M��ϫ�x�̛i�exǓ�L����'�J���\��v��%��ڻ�)�E���;���v)�)��7;J��|�{����Ց7��Gdl|����ݣv&!0n���K�r�/l�S]`Q紊T,p1Y0n�%�m؅,��C�f�z�g���S+x�ɹ�r3�c�ػ��&�`�o�V�ʬ-nW�L����2��4ˎR�X��ӂ������wEΜ������ۊK�&��C�5�_y�0�o�wHq�D�=��)���tL��ʔw�ڱW-��[d��ՇL��bӸS
ӿ'q�D��:mXڰ����9�"�j�:���>�p (D�v���|-�5We	%,��������R�)�+��g4b%��fG3�;�L���7bP��J���T6K�1ڢq���"�+3��q:-׉��tgx����v�d�'*+N8����)N�a�7�|�
��G�J\b�9�qr��9�y����Z�J�S
�d���qC�.
���\ي2��6Z�9�K�vwNC��[�y =v�����J� �x���,�W��T�9�xv�C�b͘�2�X�*�K���H��-�0K��Y��*,>3"�
��l�\f��ң��PE2�n�{9��5,�$C�W�:,:]�4T���*��8R�`�9��2�{���>���c�	1 q#L�R�gCH��<�T����q�\����8|.���s�����{*�J�pn���^�>�r�c�S���mmtF7̌^�������nѷX�At;�uD��:�v�]�ݬ�T�V�pƘy��XN;q��\#�;Q{Q�,{[�瞠k�3�b�v;J��&9��8��c����щ*�X�릥���r��:�NNë��ճQ%{[�2���np��	Ν;������v���෶���ﯯ�1�]� �{l��ԥ���uخ�`ݺ��5�k��]l�nN��.�j�ٝ�}����c�|��Ҿ��J3�6d��r,:l�k/嫰B�aI,�^b�`�s�i�T�W���q2��hٳmB�g��d���V6���{:YZ������9�����6o�iC��9]�i��S,b9��&i�/��'!��\:s�����t]0қ�ظ���I
L���1�������Z
[��Z�wS�U^*�㔙c+�Y�:��������D�)�#sZ�U,N�����î�ϕh�jѹ�Uf(0�77Q�O��ۢۗi X7d$����S��wWp�9�,r�,�i��T�X�rB�B|sp+z����(RZ���t�x�߽;��b���DI����q�D!)9�|?o�w
��;w���!�W�6qB��2��5�Ј��@��;op�æ������2z�31�nu3W��J�AtX|Y���e-u��W��9^1�oW�x��%�YL�:Ԗ�b�x��ZwNC��q�"�NQ�Saޕy���3�je(!����P�)��/u2��V75aLC<Ud}�ߥ��V+�qg���K� ��u����9n����m��t!p�d�\� ��y²�;�t��2�u��(aLӱ9J��jM��Cx�Y&&X���GK-M�H�;�9�L��Ӹ%�l��\��EdjR�猿�0�>?f����Z*ݣ�9j��t���oU3Fi�lS����W��Ep}�Iբ&���r�C�:q�r���Xu�m/�4��{��"��He�X�u��K����J`���|i�!�:|�w�f��}rxP挤G��b8�wCcN�ӲZYgp����މ��<s���&V��[5aPў����9�-˭�4ʪ���q�-��u�\�\vt�Y�Ѣ���K\�Ok�
r�8�"�ȋj�Xt����J�Z3O���S4g�:��T,e#��~}��0����%(�i$rID�C<V|��rHg�ˎq2�sķ>t�ã�����2a��&�bfe�]���U�7�b���Z��U3FȽj�󬞵�h�TS�]�U8�V2[m;�L�w7�p����ۼ�����J`4��NV>Z����r�II��a�rf{b�0^?uk@����[E
�~�)B��1d�����_=R�CFs�6M�)�9Y/k��e7m��9b��ֺWc�&^�\�q$�mSV�5�:��Cs�<�r�7��ťS+F")7���4�76����K�R�Aa񳻢�tܫH�#(�����0�����!�<;������R��,f�a=�L�`�s��elnQ�M�{�0]?Lߟp�)�v�B�T�tϜ3���SX�.�L9��wZ��y"�t����D�xv�bg�ٸ�2���f&i�^?v�Ӻ/��3���dpn���ڼ��
���`����8�����S<e�;J��%>?�ʝ공���j�ۄ9��H�   ��B���r�e���jR��8F̔�z�-p��6���Y��vz�bM�k`�>&n�����4[���%����r�n�u��4�ݝ6���f�틮	�O+��P�ͺs��6�j{#y�;�XS��ㆮ�-Ѵ��]����z�X�=]�I��88eS�\�Î3���l�WWF��ƹ����YSV,��s�N���K��OE��K�wF��;��a���i�'j?�?Q�st��S[`�6��[����GS��tT��{�Чj���{%ּ͖��ݷ6�/��yt��<W����0ex�NZ�f�=�k�
ў+���X�+��d&��EQȩ�<aϋ�{��r�g���&sFx�/uS�Ec�m3��|=�mn'���,�ws��҅X�u�غS0�f�ܒ
X/��ҋ��@$5�6�R�ۼ�9c*��RZ�X�8ٓ֡�)se�U��cjZ�!�3������emI�e��4������xÈi�N�"��̞�`�|��S4g�˙�УP{ʛ�:ʢr���;X�*;A�jz����s;���=�qu���������M�-E�֣	-��x�3Z�ے�(V�G�gut�f��]��S0�W����*֋��+�3_�辟��%�@�Pr.4h�9k��QtjѠ�ikv��7�{�LC+J�7;I�2������9���n���-���	m��U���T�9�I��T0g��o{�������9��;�J�jIyd���T���8&!��#S��3�b��ʱ����z�����T��Ym]���}��AaӋ����P���Rb�X�9.Ov�0etU~�7�ș-	eU��	X7Ѯ�l�^�Y�\��ju6La�ڌ�N���r�	���t�MN=���� �����"��p��`�x��7�S<_��Cm�WZ��m�wt�����U!�s�RR���"�PP��Ѽݫ�%��w�m�H��I[rQ�;�h�Tq{��g���fݪ�r�{����U��n^��	6�~V��ݼ�<9S�^Z���Uٵ��0�=A��l��vVޢ��0����w*�:�f��������$i����e-ʀ�w>�:ֽJ��޽�VH��c^��m����1yY�9���rwb��w����*�tQ�m�dvRR���^:Z�32��[��u:�j<@xĎ�w&�;���N�лܻ�pBp'.�7���4�%콬�R �3WB�*�m]j�A`��e7�.� dJaUy�IM�����1E����O,nԠ�>2�Cp-x�AA�d�5�釲�4��\`�����E,�(�Co�F,����tܷ|��ɍ�u���l�7*+���t��f((#�\�ח�kF����L�FN;TڵH��*2ކ�P��8Y�zի��V]��t�	f��	(�J�F݉�oYDՔU�n�0�w�췇���Z7R(K<dʷ�Z���5��O���]xӓħӅ+H�b�&�i�B��h ��6�'��,��eb�q�m�Kiy�T��(]8��zP�����P^�v��2��}:�3�e��.�e�n�;n�v���&0�S
��)E��*SR<���F�B�P�Y�o� tI@$�n
h�r@�uѦ@ -���0X(
*mTbN��	�7�2��U�
ثR��lR�y99�}z��j �m�XE1�&�7z��;�� �@^�w	�Բ��=������(Pv��L���0G��U�D��fa����q1-�Ü@v��P@��H����o����!�û�έ!��l�96����BnJV�}��i�L��Gbr�*�"Lܙ�Bt_�������7�7J�r�H]v�1B�b>�=�L��"����g�N�!��/Eq�9-S��}�E��v��{]۰x���n-A�-���nz��0U8��88�6!�;����X3N�d]*3J�I���燛��V7|w_V
xtY�knZ��r�HS�a��o��0_��u3N3�|��!�+>�E�!�+��'Ҷ[J䖃��y�:aύ��t�����Rg0f�Ԙ�2����(C����[�-$R�aN�a���V�C��1q�1-�	�2�n�5]�$5���T=� Òx�wâ�x�tnk�����e^a��8�x��U3#�=&�CFW�r{0����!�r���ݮS�n1^4m���z�x��`r�V��v0�L�McU�ų>=���w�\��\��e��;�h�+-�
3�>{;����[��g4b>s�j��4����]�IKe���J��L�����!�<Y�+x�O�\�ҺԖ�c9��|���X�C�FS�xXx���ӸsFxoT�U�:��Pє��8-<s��Z��Gl+�ӣ��E�;�rv��d��Cs��ҝL�a�����rt�7��c��$��Wr�CV��S,exw6��g����U����[_W{�}��%0�a��ܝ�@Ʈ����7�?m��\�����9dʌ� v%,1��I����$��Fwm�r��F[����^�U��臸��R�qp�n�A��,��Fc�2'�n�i�����7�;.;r���s�j�+Xxg#�q�vW!��\\�ڞ�T��� �����k�{X�f�ug�bg���qnp��n8��=M���p�<�@�;�ă�f�aC;���9k�=����u��ʧrA�M.����)�78�'b[tlkv3]���YM��KY�p���[�C�Wn�0g���Lҙ�[���1�:��8�w滥0]7}�������u}��P��G\�i�c�jJ�CFi]�RuB�sO���Pҙ���*�U,v��7e�Ð��w{��æ��9�LC+�O�u1g���!�w;��ǲ;��i)%:Ha�~��JS)��(YL��N����X���)��7����'�c����!����f�b>�=�
ш���!L>�������W~��u:�bh���#�Y�{'�U5��M]m�v��qhۘ����N���L�cm��9v{���S<v=�����n*���ϭ8&i�񳺴��.��Zcr^6B�*�-2�b>Rh����س*�+���uâ����LC��s���Ez}��|`�x�'��S܎q3�a�����!8�U�h:S�N�t�bs�2�؜�8�v')B�b0��U���b�4NG=��DevQA珝d��iLG�9�<G��b9�ʹ�2�KS�P�/;ޙEe���+
g�i�(U�G~zEҘ�i_\�J3�v��)�7EOn]��a�ą��I��[�$�>���l�� �cn#GU�'ux��oluf�^:�)B����Jш�T�T��>u�֙�)��P��FG4P��&�w�_s;u}���z�B�0g�i��A�����LE3Ir{����-S,b9:gS���V�����ot���a�t�0��7��/Vp1�t����i8G*j���rf-Z�z����N��LC9�L�
ý�ʼ�N�d��xXt���>��a����uaFiδ�҆�%�����ʧ�;�#$��Nڻ��2vn�sHa�b�2�,�W���z��3�d���X�~]Y��PB���:*�R�>I��X��e��
�q��mݞ�;8a5�QE��y�҅�����էL�s;��t�|gk�Jq��z(V���\fҞ��lN��$#���j�Þ�t�S�l��0f��I��c<q�͙�!��D�|АO��������>sz�Hg���S��;�fs���N�E��[��Ȉ�y�9#�/)T+#�{:��3N5�b���qi�<s���A���YK�����[���1��:��a��������g�M�T��^Xe�2�x�r{�3�ǎZf���C<5&�*f��g�:���gnhp�n3qn�'c����=;��ѬUn\W{YI���;�Y^�;��i���4�i֧���3N���*�#�c�r0�_�~�]���f����䍫������)�����sF"MR�B�V��9�LC+�_�q3�r�xχ3�aE��ۀ��EL:;�n>���}s��Zw�]("��i�9�4��m�-���k�2�.�<a㙵��i�#��2��"8���C�듷�X�����Q�Ҁ�iI_t���6v�,�#���`�dsEP��9����!�����`�!��Q!�T��OB��}=�}s�.�0���kbj�J�loO)��4���GM���K���yy6�λHL�^�1�6G��I��$,b�9������U�.=C�����Kr��ڊط�otQ��;�4�6ɸ���w��zf�j�n���r)H�[q�N:�WI�Ggod�W�pn��<=r�t��᫴��ݣ����E��]4�㐴9�AѠ8�<ڙIb��ΈN7, �
�W��IȻ�)g]�[�g.�጗=���luŋ��ⶊ8�W���rh,k�ә���=�8�|���eh�g�N�����Z���ؠ�b6_n����y�ܶ[#���9L<;��ui<r�k����؜�ʲ���ިVұ��։d�7���{y�0�]zwHa�8��CJb3�U2��H��Pѝ9wz�Q5OxW�W%��t�|;�!I��3O�:�Z3N����w3�;�E���Ճ�(�#��QYj�S&��T*�i��+Js6��c)8�i�q��J:��*�.qǖnm��4shn�=����L���ծt��ֹ��c��N#�gt�U�h��R��.A�ME2�,�W��Π��3N���!�;d�w�r��3,+rέ!��no~}�,aѸԐ�E(�E	�+x�����t�݅/�8�|�'�2�b>xOur1�k׭JȡVD��N������L��9����8xU2�]�x]Ҙ.��٩Ɯ+��-u��{�8�;��V13�3�CiMd�(A`�.gv.��a�k>�N��Qb.r˼�P���l�Pњs�jexo6e&i�i&ͺP��~�6�a.����<���M�(v�u<�O���'�ݦ��4u�]���qH�󥥱V�l���i]��&X�h�l�)���)T*�!�ۂ�h�9�J�;���i�e�^Wl]�/��w��<s���
��tϜ3���V9;��爦����Z��H��;�6w5wC���^�(�jnHr�A "4Ă	����$�<sv�gp���zi�!�<f�_s��w�������Z1�=k�ш��OZ���29����7��C<c������F�"��v�ua��=�wN�/����QLP���Vq�3�6~~��;�s���-�0��7+�Ł���9nλQm�4����jȻ�K�R���d��#q�N��|\���X|dݘ������h�9�֡�)ľ��ڊ��qZ�m��S�|;�i�+iߓ�.Aһ����1����a��+�q�X��e�wC8{z�3N:��,e#�iLF|��e!�5J(/;��YWgAu^%ҡ�<VG4��=]�f��7���!�?Ӂ�G>����q6��D4��b m� ���O�s���_�x���M�+++EQ��m�eh�9�����oT+Fh����:a����X/�V�n=���ޱ�r݃���\n�:�{j�=�5ڸӕu`�Өn=j�xܛ�3�S�ƣ�ͭ~~�����W�UB���W�P���b��`�;�uwEE���Y�͡�]i�;�y��<5��3x���t��9ᬗ)�͘����UNK����նޭ:a�~�;�0_���aLӹ�(Vѽ�ʆ��Yf���ܕ6X)��St{�ӺB��5v
��6j���3�1��(C�>���j-䢶Y�:s�2�g�>s{�b���0g<KNqB�b*S�m�ɥ&�ם���z��JnH����t]� a�
c��Yw��W��ERx���l#kx����Yb�r��#x�L���f�q�9�͢N	��u ��&^yN^):˺=Yy&CH�v�(J�O4mn^�Z^�6t�7v��`Wr�`�@�[�]5n�J��6�Z�J�`F[��ƭcj��6w}�P�(y߂�]i,�"�6�BxV�d�~t�Ce�:��j��r���<25:���W�U[������Aɭ�k��\�m�墱�}*)Z�x���ۚ���ƖU��l"�5��"��'u����b���������Db+O]1T�jQíЬ�� `����\���{��M�%Ӧ��E�kN5$��C:�FD8��Zk9m�FEWإ^���|�W�>W͹�fl�WW!�9Z�1����Y��	h�R��F#Y��lB�|��B����*˦�S�ʀ9+q�b�o.S�o� �0�X�=܍!wrx䀲�Őt�H�mҔ.!!�0���&�醶hN�_U���9�V^u���ш+9)�"��J��B�=���r"6��[2��}bܵqaw}t����E�+�b���%�����JDN�ܬ���Ѹ3-�t<+�}}�6�Kţ�A�������qd]���j�G���G������On�D�Ƙ��N�>c֟�y�x��U�ʍR� (K�����(*���$�t�H�{]]
�� �IQ⽵f�tk��V�);�ۮ;��$�u�*!&�샪^�p
�ǘ�=��&�
�$zN+��ηL���k�4l�s7=��Cs�u��Luu��C���<n�V��@�WO�K]�1qd8 �^�æ��n�;c�f��o@�ܨ�f��gz�Jxsi�=����j�����\\m���ک(.zV��$��{/:*����1s܉�;W\n�gu��+���u)vI�^5�/痢���nu���.ۣ��s���ĒA�ob�rsxzVk�;&�t=���u�<z�����W��<uĲZ����^�uc�l�����J^qs��.N�痳ہ���S\[�Tj�͵zQ\�w#�� �e�㖨����������Kǆ��qGmAԋ\�÷]�p����7V�JTe�����5W���^R���g�B8�94�d���f�n�!x�ضR��Vx�vf��-hǬ�`V�ȗ#s��s�J	ى�>y�v���h�b9}���񴛦�z�q�wf���6$i8@�h{M�n[z+i.���xl�7Z.4n�KWe%s�Wp�j�uE�g���=X�-Xy.����.6�#�ݙ����V��`	�u�N����ix壂9�����h9wv���Oo)�`�Nt�\&�=O��E�vI��������q��i�=q��Uo>.3<�X���v��n�ݝζE�i�H���)�u\.��s���W;g�Zܖڽvf��Z�q�λo[1�F�n���^�q�c7�Ϯ֘�n������N]Ɠĭ�����ݰl��&�5ř;]%y�Zv��ʝu\4n9�١5δ`ה��C�[pK�=mr]]v.q�����p���`�<�U��y7�g����2�jhӑ݆�h���goU1��Rg�P���b�f�x�<
�n۴xN������ջu�����f��D]�$�3m��\]xz{n�m]��N��둌���x��/����\Xy��^kqؐ�]��]>�K�ne����p��,k�2�sk������5�a7l�:�����N��Z�]3Oa��|!��ֱ��$��Q�m��qZ�<��u�ds�)�us5tƼr`g9;D�����=�l��:�������}���c���C����;U�\N:�n��m���rЪ���8�p�<t��>W����\�<�w윜s��K��۷Wn1�&j�ӣk��l�mqu6wu���r�����9�^��[�㶜�^��quݖ�aF� �lcg�Ѡ�.:�-;����u�݂�j��8⧷�G�879۶��C���T �jz+��b9�v�����"���[��>
��է�<t��mgpM9y��\�v:�r�oW��\(5r�Y�)j��#m"�\��cw]v����*VO7l95�97�'-p��^��[q��X�8��/�D��I`;x7T,�ځ�9\��s�>QJU�Ԙ�c+N�:���L���L:~�� �$���"�K�����Φh�i��j�xv���9<Y����|r���+eq�o{��y����^sqAg�i�L��-9Y�X�Tq{���q�E}�(�QP�(���,:~��;�<a�>juT���{�e#/�8�XS>2f�lm�\�H�A�N�a�����0b+�RR���9����ڻ�)��N*�+F�rH�k�n�ة۷��<�n��۝��=��ՕG�=�"[0�WkVp�7j���ui��a��^$�-B�3H��2�f�ι;9�0�t�H�sХ��N�L9�{};���cR&��h86�Wǁ��8���y�k<p���,�Nbg0f���U�|�KP��٫��Ԏ��!�ػ�9�F��u2�g�3fR�,b)�ى�g4ٻ��Xt���+cdRքE\�J�Hg��+¦`�q�ٽPC+�[�i��4�s֡Hb+骯��_{�2�������ў)���&�iCJg��^�4b#��T�1��;+�p���m9�W[K�9��<ܺ�����`�ې��q��F�d9���3 ����u1�w$�(Y�i��oT+Fx��qq�1ߔ���sL��!�QD�a-]ҋ;�N��a�竰U�KP�����f�gK���9҅|qӸ(a�7]�����v���mr	�J	0bQp�yk���/��	E���&�_�W�����]Ӕ�è�����Ɖ-�ʺ��9�����+H�N(#���Qz�+F#瓾;�<a�~��x--��7d�wH2�L�oS0�x��tT�C<vHxU�0�͝��t��C�6ވ|��Z<v����v�{Q��
s�x�LOi��=$��.(*ƨ�)m��݄�Q�{��a��9Jc��+9��I��M����J�z"l�,U�`�ء���h��2�Wq���Zu��ќ��wu�E����Ԩ�y]˳3;K����jLP����mCJg�og9��-S,b9�u'n��;k��\�NY�<`�=�k��v�B��V|�VTʯ�Q�.��Y�^ˣ���=�q�zi���ؘ(C���w�_��St�7P�$�19��9��tX|?��]Èb;�IJ��4��(`��N�B���̧��k�2��%��U���#�Xx�<쐗\�рbsU�۴����E�9ܺe%�^8�P��㎞�Ɲ._��t��^��dsD�)�����S��SZ2I�
���:aH�i�(X�G�M4�<v')2�gEg���iL>j��q�ʬbp	wX(h�i���)��6Z�,b%�����9swӸS�WA���ʲ�Y���q33�|�oT)�ӗ���ܒ	�3�v))��{2�+k���M��Z.��a��m�ӟ8��CFR͘�g�'��)xM7�RD�l�QTN�1
5�	F�#g����q16�r��v3V��q�;������bk�^\n���N��\5ŗ
m�`�k�竊1#t�ݞꮨ2ړr���\on��=��4n�k���is���&Uс��&[���4ru�0�q�sÎP�v��ncư����o ��v��^9�On��7	tAt�v]��ꮲ[����*;��mF�+�U���M�r�]v^�y����m��ⶒ��dwE�nL[:�ܒ��wIv��;��"m��������ŵ1ʵCe�K��:�7g�[j��FT��9j��5U�v޻�:i���)3s�s�
L�Zr�9�4�RN�!��)���t�p�7Y��exǏ�PÌ�ߓ�(R�����0�e����x��q���u�9���S<w ���RnR�`��{�&!��s�)33L��gn^v��KPܫ�(a�2�og4񇅝���S+�βz�4�"\��X�:ի�/U-E�P��uaL:q�٧Y�+F���x�{.�)ӭ�a�i�
�4���Z�mB�8(Z�αtWl�m�3[���F�]��Z�+�jٗ�Y�/M Yd@�6���tÝ���!L�L��C�1:�-S4g�|�w�K��=OYP���}��0�w7�p�Ɓ���I#R84��b@��>xK���;��a�����9���9�Z}����ݬ{���[B*K��]Ӕ���c)�I�2�E��g��7b��35}�����C������"��֠�qII�S<4��(s�3_�V0��[P?&���rV���ق��>MN�i�x�RZ�X�$Փ;�X�*L��2�q��u��.�ͭq�S����������:˹�]j㵢6^.-��cS�1��1��r��خW]��u2�b͘�����UAG3�7�Ϻ2�r�LG�&S�];�X;X>F����x�����}�0�݂��杊AB�b>y���4f�N��/��R;c�.�:aә����K��}��S��@� l��5,��Eu��X��
�K��hև�4�a���w�~>f��S�oނm�()`�嶮���y�pP�br�9c܎R�X�Ҿy�;����z58�V�c���Hs8�t�Z1�l��X�T��(YX.���>�E���1MK��$j�I�4]s�����L��wWZ�u��E��In!jr�B� ;S-�4�wt��s�
U�r�PC+�L�L�+�w5w</�w�ݭ4Y,��D,ĳ���V<$�r��9��{ �f�����*��ֆ4U��xx�h:����t�|<�j�Na���4i��q�g�v���)��_ݝ�$�v�e�ҋ����9L<9�pT�H��^��0<PmW���^7��[�r*=����	�À�i�f���~<s�:�[��JBګmB����
�ݝ���c��(`�xhsm1��II�F7������j7b�j�v1Ì��nؗ�p�/F�8�����48�ϋR��.������p����!��w��S��8����O]&V�C�ݝ\��B�7�nY!ImEr��<aΗ�o���g�nwD�!�:��Ҧ!��_�i�)������m�V:7��*Sߔ��Hf�2Hg!c4�㓴�9�;�ڻ�E����ȜG�r�,�;��P�Dy<*b�u��L�����)C3ĵ!Jc����˼���w������)�ي3�9�qC
f�Ԩ&r�!�6Z�h�*����{����K���A�¹nm1�p4�NB�m۩q�	����d@�FКyS����f&v{p'���JV�5��v\�H&����*���Q&w Z�2���on٭&�����<I�Sb��z�εð8�6��U�.�U��If�l�"1�ڍ�mrj.z�x�n�.�6�..8����qL^wQZzۛc�Wq�n��=������I�6f�;<t����\�쬒s��p���+��q]���Ӻ{5���5kU��.=���f�d":̣�g��gbw'm�[�;g�u��:6^޺�I�mt��N���8it���,ex�?=j�1E:�V3JϜ�e1�]iˤ��2�,;�e��v����fe("��ړ2�f�)4U�<�i�2��%AB�3Ir�X�KYk�����?n���<1��i�g<g�N�"��&�T)|~��v�#`KY]R��)��;���f�;�IJq�d�uB�g������x[��q��Ei(7e��C
ex���)��E�sF"<�1G1ɶ��+Æwj�K2����v�m;�Z�v�u`kˉ�ˆ'n��]�J�틴4&:�g�>�t�qud��m����x�6v�*�#��`��3Jv���>�4Pҙ�HR�`Qvw�w��Wp�L<b�ݽZ,��� �^=�/>bエ8��IsH �8��1�<s&�k��t��ڻ��a�����������X(�l�w�,�!����qC
eiߓ�("����8�h���P��s.��s�}�:��,��C�{wE�!�<f]�Reh�6E�\��Ee�:��9�H�C�\�K�Ԏ�gt������ե`�����!���u�2���;�9����P-�J�ʘ0e#q d��7K���Ȭ9�`I�j�AF�`��T�+4���(aҙ��y�Fx��S���9�It�e3��纡�0�V��6�-@p�K_V�0]~{:��V�Iz(a�x���&R��ش�0�Q~�H�A�E*���Jg4sf��>��J�[ʼ6m�myf�]��3�Vc�\����u�vc��Ν֭���:fXi�����YV"���+�"c`	�%[�����8X��q��@�v��_�n�ؔ7BE�8f����e`�VyҤ�"E�^��Wn#R�ЗW]��+!�J��wg��7�_<�B��V�˷'��b�4���L�]�Z�gBর��]�4�b�[�agg	�8���U�E<Q]�^�W�F�V�T�3�'LjJ�l��6������`U�b�Ӯ��
v�/����N��칃�{�il��[�̖���h�	I,��esK*�v�3I�u���'k��͞4.���0Y�\-D��!�̳Wv����Vn�z�&T̻��ۈ:�a��r�uKk����cѶvU�Ϋ�f!a�s%�d�B�8�r#v���E�v�v��&"I�I�1f)�X �L*%�)'GPPM{EE��XT�W�&�j��eS���)�דUF�w1&\1��캍��x�� &H���B65�X*]��Х}��"t��\R˨�Wg^�d�,�MZ!�fV居���Ur9D e=�{f��m�u1�	�1ܰP��ߥX���cb����'Gd�.f_�����ݫZ&˓�h�-�!$�v�B��`�u��*�Ǌ�Nv�es�����$��Kt�
���ϯ��1�$�v"F�Vu�b�̛E5�9nm�YE ꙍ]X^�,�SZ�����4�y|�;O��^���kbX�%��q"�#�/~�ë�����ٽ�����߭�ʩG�ؙ���֙Z1�9�\�⻒T;�0燽��t�æMg�17\l�2�yۼ�P�G~�)T�q�s0ex�d�Pӌ����(V�C�R�~��Y�ؼ�'vҬ[�(5�V�Ýq=��E'�f����)�6[s�sahz-�^f$T0b*<��#���f����C<u��
��R+�|w���%�V8�Z����绫�.��4L�3F�d]�4g�v��B�sO�\QF=UY9v',�X|~˿N�+F#>sz�g�g�oS���ӸS�|n��~��-�
Ky�0Gq��\fҺ���aL�v))�b�ŧT袨�F�5D����C���8����43���
X�eD-����a��"��h�G�M+Jg������ï��ҘxV,Y��w�Ψ�}�܋vՎ�E;:�S=:w^skR�q�^�]�KqҦ��(((�v�ȝ���ӟ�~V��S4�}%&si؜�P������<`�<�=M�VG[$��,�4�:��
ў>y=h)�1-�
3�Ϝަ"�����;�]�s+3�f_s.�9�<vHxU�I=��Ӯl��8�u�-B�f���k���D� ����0�N��]�sO�N�PҘ��=�`�I�TΜ���0|�P����gp����q2�1��ΨR�Zr�r3J�nj�Þ)P�����"�Ü���x:�<Cү ��
Q(*X��w�kjڬj�EZ��ըONZ��[����q�x�;E�aֶ���@�ݻ�{M���2�y�����aOZ�)R��G��Gn1�3ۛE;.;�l�\��:���uu���Y�<v�y�l��������|���s�N��(����ݎ�\&qu��Ǹ���mtۮ��Eu��.���q�1���Fݬ�5��[��-��ë��T֢v&+�L��$�K�ڸM+%�7M:��]�a��APɚ��ӧ�����Y{\ޣӴi�GE�a���qkj�j�'���Z����sK�5_��
g�y;�&sxv��UZW�/E�<`�~ۿ��0�b�{,$R�Q���gS)�Xږ�3�e�8�c9�T�)���P�FBM��rV��V2�9WV���?N������8�����12�b�~�_N���m���KGe]Ҙs���f�jK�L��[��e"��ػ�0^3n������*r��!�#�Ii�c4�㕜���Mgd�0�����}����{�Z��u�[��<�m��5<%���v���*���y�K��磊��W3���$G&ٳ���~��H�j��#���Lє�nwD�q�����0���ƻ��VYT��J�a�~��]��@��0p��\��V�AE�nc[IM�D8���;��x���iS+F"L�t�1l���e�JJ�b��w
`�~˿N��F8��U��Y�S��C<W~��(#t����-��X�cn�N��aὛ��ў:��T�H��IJ2��0ӺS�|n{���Pv���u��P����R�4b*<�L�g�k��t�0����~LS����Á�������{uN��v�]q��/5��'�ػwk)6h��w�tw��!�9��0ei��R�b͘�Va�w�}g4��<֧��Xª�{�̤�)��{�:��3��'�h�K��UH���S0exp��3�^e�Z�+%���!�>7}���*a����ϛ��鴑%A�4U�3��X(k�9�<u��CI \m�x��~]��<\���X|fxGCk�RVX�nIJwS�I��c<s�|(h�G�/ZeiLCޟ �~��y�KD�`4!p�!�<S�OZf�;�8R��%������͵Lў9�����Y3�/3�h6���0૮ɦ��u���W\��8�u�4��6wn���\�(7�I�f��$2�|��+Jg��S��Z3�H�P-!��ݻ��Ý?M���$
�>����u3
b1��8�x�攩�3�"r�L���[�i��4��>���v���N�a�}uæ�.�4g4u3f(YLG\�i����M5�!�E� �vέ)�N_پ}b^2�����3�~zAB��r�ހt�I�'�V����w66����U�((���[��w�Zt�����ƾVG�D|;y�3�}6h��3N���g0f���_V���3+�����g��n;?����k��yQ\�F��mY����s���W�a+���+4^^6WsY��4��/ΦR�&�r3�uӞ��3���P��&�n���3�w2�9��$B�x�X�&`����q�6d��V�D{�Ew*uTAIc���S�f�ϸSt�M�f�9z&q�z��3�6�yH��RT܃)k�0_7�T,��l�
��v� ���;]����X][$Q؇�!��N�1'7��ў>y=j������Lÿ�E�)�<r����l�� 1��똈����V�XѠ�͝U�j�n�m��H�~w�㜫��Mq�Yvm����c����W��b��ֻs��u������o�擰�1�@��p�!#�@֮)��z�9��a��N��\]Ws4�r�
;&�]�c��N�rC��6Q�O[�����u㗎ܯk��e|hڕB{�3Xz��y�R�۬����3ѤP�v\��F��'\��%u�I��]&;��g��S�qς�|�����q�C���|���e���F���nƣ�
�HR�C��i��ю��/,m���u�<��'kb�2�Ơ{A��t~�����-K�!�4��%�X�i�6Z�.Su�NC��P��+ �;y�gUCFiƌ��,exs6b��b>�=��ш�������d�U��ڪ*�Y-�p��|~�i�xX|d{13�f�� �3N|�e�h���xP �kpu��l�t�0�qovw
��>xOuq�1^��g�N�tX|~�t4#V uU+#$�wNx����U�w���>�R�9�û����,��m�',�N����c�u��Ӡ`��u�DW���:�um���X�{6�x���1W����Ja�MN҆�珜]�1��&s#�_l�����7ɽd�h�X�v��:`�2w6��B��9I��9�\۴5lMb��M���0F��lV0���"�|�^뭝L��{+E�!�VF�&`�|U��㕫���e�Z��E���}��9�ٛ-S4ei_=&�CFW��ON��t�۲/%
A����:g�gJ�ұ���xϝM�b)�7~}Ôã��	�E���%�S0b9&l�H�:���q�c���U���v{��ш���+��;]à0tޫ�qw��nn��Iۜń�hbJ�3%n�fd�-�z�:jb�����29����7��C<u�{��F0��wn��t�w[�HQ�X���ڜ ���:���D�oT��)��N�9�r���Aa��lzD!�Y,��M����8A���+��b���{zݧ��b�)�*�F�5���8g[�kr��[c�� s�� ��q	8�=ۯN�C�|l�転�7i��4B'dt��}��W�<Wbr�,gӛ��xv�'S9c4�/v�AG>��_Z�Z-"�$��`�n�l���S���x��p�Cx��M)A��Xw�d�U9+,UKa
�x��60u��e��G0�a�F#���kn��Id�9Ur8�.��a�}���ELў8�I��2�Ǐ�PÌ��Z#��DU-��F펝�xå��J\���w-3�9�>juA���k�r�|d�~m��+mq���2�x�[��A�ٸ���F�,0�λ���!�����m��sx�'N�yjS+��T�Pҙ��ي���~�ZSp���i1
3� ��	�� �[TUF��DUsd�HQI�ڀ����V�w�i�)��\��%mG,�H���Wt�0�s�3�N�3Jw'�Cql�P�s�}������r7
j<ӝ�5�]���vgM�p+��zŽ��Y]��"ZH���[�T^w�h��I��c4��T�Pѕ��E8�29�e`��2��,��lECr�Qa���q��)�<?�uS4�NZ�0f�oe���2�~X���J����Ҙ/��]��3F�W��Z1�z��_[���s��7���h����-�ҋ�N��g0g��oiS0g�9�����_۾;���w�-���G��+i��s�)�3J�OoiCJeh�f�L����8�xʧR|fe�%u33%�,��^�F�'��CQ�&6�ՓH's7]F9��>.u��ߤ�m�!�tVf*4�n�݋����t6�J9DҶ{��JK+��W�r��Rvu�Ŏ���_}��R�	�LcC+	˗r*8���J&���;�i�JI�
�� ��m�R�q�vV�r;�k�<M抝��Grq�h��������(��SM4�8�܋���w��W5��nE�u�j&�
���E��x��zsIi��i:!R�q.5.*�74���@h{n���j�(T]2XTAftY"��<���a���{b��i���u���F/�$X�v;����(SyGm*�j���1��U�=��]֕	�a��&��)�52�콪�D�(��A�&ߙ��Z����u���N���7�a2e��3WR��V�,A���e�.�Uل�A[hf��*ǘ��׀��V���z�ud%ҝJ��CT��P�F��Qk�V�(�Tu2�>��:!�R��^Rl��
"j&=Ĳ�^*S}�K��q0Z6H��YL�Yn"�����]�]�T)�ю��wr���3l�*-���Ĥ2�Jj��E�
Q��oPX�7m���{vΙ��#LSzc��d|v�/���+%�\� ]�Q�P5k�N�;"X̓,�׻=qЀ��nƺ��ܛ�!t��J�Z(�(��h�[]M+˗�
ݭۨ���,R �*+���^�g4��7V���Ef�mn���A��A�|�ڌJ�+�γ������gj��ě���oE��X{����D�t=�o� :���kn�s��cp$�wc�v��X�z����W�^۫��*���c��OZ1�y�mrʱ;�wu]b������.GoM�f�L o=cevvƧ^����ωR�KE5��52�m�ţm\��j�J��_
�q�����e�m�g�A��tט�t�d�ۛ���l]=�8�;/��j�������=)y8x�nzm����w��@����n8��B�{�p��9�6(��i�=^6��v���4v�;��I
���n;x��ac��c��8=��)�\z7K�Ag[΢�'\��tQ�o`������[��5Ϸ���7	j"���-]��8�=������쵶;"u"^˹|"��۷u�m�7n���6���g%��F�&��.��v�8���bKc�{x	p����{ZZ:6��v�k��%�K�����Tj��:�.5g5��2P�gUq�0���`�LLv���ͩ&E9��藻G�v=���.zT��ŀD�nOlcL�fڷ�DY�W�I�n^o[��pN�n��蛶T��P�30>ճ�3Q�u���9o)̑�f�́����Om5������\YIkvqn8��^��F��J�a�;��vusd�-u"����4�Möl�K���)5G�s�Lc����]�s����:����9Vݯu�Y���wT���f`�2.A�v{<\�'�=�����ʼ��Q�����`��%a�kb�e�n�x�k[������h3r�r��@tq�>[�um�/nH�;�cĆ���T�g��?T'Ǿ���q�)��9����Zۀ������G�N��7����CBu۞�Mc��qj�N��.���Jy��5nCE׈+�p��!烵�O.��q\S��U9�.�@�4(ڎ�9%8����F��e+�88d,n)pp֬n��W�6�u�Ǝg��nN�i{F:VOl]]V{k�m>^����կ����NM�On�.z�Ҷ
�ư{#��v��i�J9�t��s|��������v箨b�^��Y�%k�Jb�'�|}�� x;��]�@�̊{�=�y{��\TQrԷ-<��Bљti4#�����)UuW9QR�
�Du�z�a�=�Ѫ��eI��$�[�S�K��L㴃�];���p6K�7[5���z��VN�s�h�@n�kOhť$rn�Ǔ��[�S����m��n�*i����0۴r��q]7�A\�78��3��v�Ho\ ��r��͞�Fs4l0�ס�Gn���fу]�l�����u�K��g�c^�1�v	�+5u�Y9x��s����/\�;z��Y�]���`�&k�;c��I��K����q�akZ4kN�S�FPl�:�Z��������ױ�Ng{�~��|i��������R;�I�8�;��P��NV����VU�/�p�7�nT[%;�0��o��E����v�2�f�:�-S4g�4d��c+�n�kQ)B��6��Oç���+F#&�r3�e�8�e2�9���Xxw7k�:&�w��ae�Ðbٸ��3N5�be���PG�:]��0�y�W�9
�kp�w���v�bb�1㖡�3�NnR���x�L���q�QF]�����V�h�q�������h=F���kOUD�u!��Οn�\�5�v�):T��ީ��q�;�)ѽ��O|,�y��Q`�~[����WUQV�#n^wO��}��&@$$;c�2A7[�+�Tܱ���㉍��9�؇N�S]N��3�\�i0(�8�q1~0�}�q�`�#�8&`���p���f�x(���Y+]�t������"��II�3�9�b���;��T���.��pnh�V4 勫Ox�9��h�D����q��s֙Hb:\�w�C{�j�vF���x�c9�'PPE3L���`�d����|,�ͽҘ/4��V"�Z��������!S�Qu�� h:�.�8i�Yy�rn�uf��`7`�����b�3FȽi������Y"�ZC|os|w
,<l׿ZՖAЭ:۾�uS+F"I�T�3ND�h��+F��L�S<w�=��C_2���j!�Ƨm�o4�
��k�C|d����O� 8 !��	��`i����퍶:؂���2§p/��}ʉϓ�=}�@WK;"�����T0f��M���Y-R�V��p������ӌ�,��
��v')2�"�����gnBk%j"r���đz�3�b���X�q�͘�cO�w�x�?j��n9a-Zt��m�,l�К��.��d��{�-���`��x���8��t�d�E#��BJwL>)>p�Cx��{z��sH練��f�w6�S����VېRYj���i�L���[�:������+F!�/Z�4b+�z@,+�u�}��K�Φ!�FG4L�&�3�3÷��b�u��(`��/�:j�5`8:�-]�tXx{���0�w7��S���ZwJ,8��|��!IV��F�lV�i(��$��i��Z���@0C����$D��-��t�ã����ٲ�9,U*�}Ôæ�ߎ�:1�9�Lѕ��e�f��:��#��Z�jq�D8P�����Ys��EL����l�uÖ�n&q���F�G��6dmZ����΂ҘxO{���0�G6n(aL���Φr�!�6Z�X�sb�o*���[p����߭3N1�oS)ҳ�7��C<V}%x�0��ʞhV����-�+_pҙ�M����#�Ij�c4�\r�!����^������!���ʛG/r���2���O$T0b+>��3�3�pPE3�7;���I��}[WC�v��RYՇL:q�sy�!�雪b�YLӹ$*�i���XT0f���c�:�\��5RET�]ju3���WV&����Qs(�"��& 5��E�v����nU�Tq�b�n��@SmkvD'ngڨ�Qh��je�n�4����S&f�4�n³�m�@r�`
��F�6�������\v*�=�c�v��	���gi�[,�8�3yI98l�qwWq�Ks��� c��85t�$�X�O�:错'��<SاY#����I���lhy�������s�mA��gP�%][U�p��ಌ�����Ƹ����:����/�aɶ�zY����-v��p�..�wl]F���5]�{F�3��M�Zl�X�wO\r�����x��|Y#%g��YL�.l�U�D��N�)�����)���=�mc���˳��]���!�ٽP�3�{�:������`�#�E)�7[7�1�%q�$B+��3� ����҆��}"�T4�-�	��>��PX�i0��Ke@T�{�0WZ��e�杓giB�b;�Ψsi�������׫lMZPvZ�\���^;���aLѽ�P���ۋ�B�"���A�>�,�{eҰ����۪�uF\Q)�^������ɩ��iX��u�x�8n��[vyb�j�3
g�rmҨV��'|*fG1��(!��))Af�MW�
��fw���b��wE<n�]��|�B�` x���Du�skTkmU6����Nn��s��yb"�!"4��(&��! n�aY>_q|h�h���L���sf(r�t����I]��K*�Z����_�7��exi��1g��nReh���k�0釅�uH?��Fӣm�_t����R���ι��`��d�!��b���.�\�M��X�p��ᙔ�ZS<}n{�����o9��&X�x�{8��1S+��ڸ��X�b�pZ��&b�n�Ɠ������78�x���\��m���yj�WD����]��4�RZ�X�8�9�2�˒��g��͘�V1�(�}�q��T���Ha�<�l�0�Ƚ�Sӛ���3�C�j��x�ڷ����-Cd�7+�0_3�;�Na��o�wE���>�� HQ���ְ���cDs+�h���ٶ��hh�H@��5�gH��}t�����k�xß0��)S*vVW��0PE3�H�U2�g����LC<s>sz��W���,��|2szUٝ���Q�EN詇�s=�z��xN�)B�ei��)�1�N�q�߅���clV����s��GX��K�fu�N�v��<;�WI������K;f�-Q�Kc�9_V��㟱]�wO.���,���Ze!�V<�aP��+�{�e#�؇,�t���ܚw)�w�%*�!�|��CFV��lŇ���7����k�

�h���3ë�1B�b�b¡cRd��`�]/��>��a�cqϕq�J��]�i3�3�[��b9���(h��zwN��O�`$!#�B@�;\�T�EM�T4DT�U��E�h")b-�Ժ8����߯pP�x_�k됋�aY��)ub��X�+���2�4��PE3��/uC�1��b9�"�{��A�n��W�G]m���m��6<�1lY�u�V���q[�u�vڈ��a�W�!��wsy�!�<l�転���;K�����l��>���*z���咝ҋ;�.��a�3z��Lє���OZf��u͖�VS�3[�U��R�[�Y�0�W3|��!�)���iL�4�7���x�fk��?Lء#o��p�J��ш㷳�Ӹ�8�1��J�uw_y�0�Y�.�6*Ԯ�e��^fu2�ei�5:��g��d9�4�)N������!I�2��QU_�b�|˃��W6���N671��ѭ[h�i-���p�%�s[�36�9�����]�8��*& �������k�n�K̾�l������&�s`�݀��;dT���\D���ی!v�ǋ����h�Pv{���-V��MeX�l���P�z�@`�*r�ص��2�o
�z���e�:�ڡ�7���˷�j�#�o<N���mU܏����\p��M��ܖ�����<76.�8#�^����v�;Q{`7t���N:����un�z���G^��vt�y�s�RY�������vE��Kv��W���&2F)�8�y��q��uż3�X�4\qf4���#=:2�#���ݳ�ÿ��.��ˑ_!c<S��3�6Om�h��v�m�(��H�l�]X.�|Ks¦`�Ew>pL���6�҅"��4x��4ѿ
(�B��Yir1�͔��8�6n(aLӿ=�]Ý0񓻵ui����D2q�T��w�s-B�R>�{�q�ϱ�2��_��`�ߤ�J�R��.t%U���H��:,<=���Su͖�2�YrAB�W�xI�9��K*:�;+�6Ig$v�[Ij��]��X��� ���D�݊�l�Q��WU��p��P�M�꧴^0�}y�O�)����q|��WƟ&�E`�.�@Z�*�2'%�V��3�o�v/�C�1�k����5\ص��1KEM�N�5��G#��r%��E�52bCi��8>4ܜ�tP~������w5k��˛۷>�I�5��Ya"!���o]L��o=�4�Z��\ǯ���Oو�t���U��+Y�=s.ŷ67�D��ږ�jM�oI(�v�Ҭ,�:ܶ��}�.n��3��o�۞����7�غs�{�x�a�i�IP;�j��k��'=��ݮՈ�p�gT�V�d�S�c��T6U!a,f�����}�u_<M��4?���z���֛|�x3�u�Y[C��c�ui�s��n�y�[3�v�w&�˙���?��^�z�貜O��W��e���o��o�a�����5K�qR۫�%�wN���tԄ^�l4��l��+�:=a#�8q��x;h<�.�%u����	4h�Kќ�K���j P.�:���2��bކ.�ήz)�w7�)J�hނ�e�W}��ƀ��z�E* nU�-8Z�V����/]�ܼv��@�g.����֡;Sl�-��5p��ɅC�WY�g�@鹷���٬y�s�`�q;YYa���JeR4dig6���5�#)���Ü�yyn��j�!p�����G��wl�ԯDU�+�H�X�8��n
s��ٶ�DL�ϱ�`��8�N勗~��q�xH���2�W���~/���,Ky�/����&�Qm��zI�[zu��WD���r!�vG�b8�XAd�k�h딷t_4���/fS�)�R��V�ۿ[��Ts���hU�V�v�Զ�ø��6dt.�
mR�00�X�)�t�UbnSLfJ� $|�	n䥯)��F
@WJ���t�j�H6�!
�暎�Wj�E�ő��H��M�<w�M۰��E$�N�XG%���T�Ҡ�ټ�Pbţ���
����ˮ�Q�)���X �P��k#�D��jt4��{�;bw:�D|8,m�+�)K���=�reuu�{���)G/yq����NX h���!ŗ-$����p=fS҃��LTnD'Z�q�*,�ѧ6�t�B��w���K�vܑ`Ǌ�c��]X�;��.����S�T;X����~I���kך�\I9�G[4�TTM$WV��yj�*"��*���PDDsj9�ɨ��������I�Á���ƙs�n�f��q�<�,���WC�]�Lxy�/�=���Q|��d����m���wnY6�H���ݒ�Go^_�޼����jZ>_i3�Q�O�͗���	��gK�ţ]��q��n*}�m=z+�J�r�k�K;n��'�e5ݭ�)�(��|�o��ǧ4w����_}�wp_Z�z|�OM:h6Z��=�]�r�����nL~.9ϻ�x�	m�PaQyAR�m�v���oL��r��?{���?nw�����AH�����%A'�ǟ�޽k7�?>�{�u�Ҁ�4cTi�/(*��m7��A��y��%]C���R�Uu�B�\�UTP�O�~�忟�����Q�E`�*�i$X׳_?�}��O��5N����R�-���?4+���7Zn17Ubd�22���z�ەOFz�8���s���c��s۝0��$,)U��S^Y�]{{e׷2~����ߝ٧��~w�#&�B�%���&}*Kh�)S>Ϣ�'Z��;����dhiH��+e��3	����^wO}��-��{�����E[ *I���;����}�읉��O'~��*u�������t |�ܪ^2�E�s���_��8��d���W��ǿ0�^�N����
��A��kZ�cEb�
�\��b'cSBrլE1D�U��T�*bf�泂&���˕�q��է�E������Nў%9�v�����l%oW��u�=l:�[Y�ꗁu��+a��^�v�7ku�C�P5�÷x�]�.۫�����a{oD�Q��K�v���W�GU�
�\��Z��K�b5*��k<���i��Ag��OjӍ9:�;��hK�ӼZ��ح�j<1k�\���X�B��nd�;���n��{b���{<0q�v�j
6�����Ŭ7;��<���vަ]��\<M��Zע�6��j�br��+[A+�Z��3?��f7;�;�N��k�ɣ_g�d���w���a��ZK&?|ѓ�}����{n�����ۙ��Ym���Q9-����;���Z%��s�Q�D�)��������J�%�n{?}7��ߖ]���[;��7���93^ʫV�2���/-���>�TO��.���7��Ɖ�g��&6E5I,(���Q�"l�:
��9@�;<��j�pc�Y���abc�{wJ��V���y���[���sE���r�Y��>����w��ݮ���伕�7k����7���M�! �p�8!*�sEU��2\��F�USCUSLQl��#c�D�@r1͈(MTS��=�Zڟ�Ŷ3{�\��.?���T^��N8
���nj�����ٷ=�{�k�~7�7��nŌ��:�V�Pw/2w�ܹm�[�w����^>�ٟxS'�j�XI(�SrgI������ͻ3�f���盵c�ם{,DCu�4��η+;��ħ;��{Y1�+Sۖ�`��|�;�xθz�y�,ٌ~���y-��o%��K��.c��ٽ��z�����n*mΛj���~�{s#���~���7>9���H)"�0�Gk����빺��ݾ���W�A�TE45F&�
�����Jb
�����QAESQ-DRQTUm��m	����! �I�����2�~.������ȡ�R6H�^m�&2_ȹ%8��$�ߔ�R\�_9��ކ��iA&����}����X�k�&lٙ37�/�cYݮ�T7eߞ��jӱR�r;t�p�������+�:'�UG�7W"��;(��B[]?n_��Wb�}.i���c��g��}
�C
db�N;�kg����^��������|�r�˫���&�F��2���$���J���ds�Kx��߰�ʝnj�b}#��'%Z�{��nw0���~��{�����k�L�X4G D�˜�s�7Qmˁ��4SE��U:�X9��4UDmZ�g�
�&�8УbL�m����<��ov)5Z7j���I%�.z?�y���7ܝ���i�ȷ%}�N�i����)؋<;,Ϊպ�p�ɨgFE���p)A�&n�q�+�vtmk��PM[�߅;���jJ�-���4��e���r�9,��R7k��3^��˔�7<eǦO�׹�s�щ��hX;Z���s�/E%D��j�L�|�u��ur^?��q=C탔c��G+���g�e�~�橏��9�~S>u	m[��]���J+-jJ���l�Z�?;��w�I�u���=�կ��`��_! $.Wlh���h�m�E��l��LV�9QPű�"�(�����h� ��8CH c9մ=���Lۛ'kWS��z<C���;�9f��%r��&ɞG�$J0�KN�����[�1k�������H@�m��Cɬ���u�on��\�:�k��0۱��d8F{v��F�[����O47���p�&:�n̽��z:�ڌP=�g]�y��/c�����c��2yMעkp�}E&�l��KwT���0����nf7G9i��ۚ���u]n:��V�Y7��r=cn���c�����ݳvNR8�뱕�mi��[�݂�f�e���S��W�H���sF㛪��-XN���������ǟ_5�:�m�u}ӻz���t�!:-��,l������.w�m��z�.L}�fWв���Y�'k��ܱ��l���ޛ3&f�~��n���r��ԝQ�U���ڙ�߰����ܓ'~_g�dǯ���w�]����KU�Yn�3.��_�nM���q����f���>��{+�6U4������WO:�n��wX��]$�͓ur]d�ks�=�`�Â�͊���O��<i��2g���r�9r�E�Bb�W,W�P��n{3o�Ϡ~*�j���sp�~j ��յ�K��MF�1�蚵����� ���Q�\ب���(��5L�"�M��o:����־��|��n�+��2H�r�:l����ز���l�O�6f���[_ۗڛ�7m�AS�\���ş�?�]���\�־��f���~ޚ;`��PM9k�����>�f[����R4��)��g�������{�7h&=r��֜GE�e�@�;{b��c�oi����'	!s�I=i��_w��ٻ��~��G��㯻�k��+��>
�D��d�[c^ޝ��:�ݝ6~��wv��c�������3U㖨�
+e�טO۫g���3Q� |zb��b�-�LM33��LC��ڊ(m(��уA�.�f���:��*
(m���RPDRQ��9Et��:�{r��{=*fɯH]��*�6��I��͋7�Ϭ.�p��7�-6f�u������5[eU�+q��1Ƌ�T�����\��,���K��kU�r@((�"��M5*r��S��� v���z�V����X��js��i�eC�K/Ĥ��M�����.]�o|9lֻ�s����۷��(�v4r�8���Mϯ�m�\Ǔ髵3��Ks�+��O���l�K��i���S�t[���mg�}c�ط������uK�^m�h����V4��L��=$����/��9�ĵ��ULlc��T�N&��"�y��PQ\�(���` ���#��C\ƚi�N�"J������K6p�%�[�t��o�gn�A�"v�ޕy˼˩�m�VH��s7�>���x�����߈І�9���r1�V���m=	�t�g֝�nuc�z�kUۮ����!cn�H��r�>8;h��f�����n����.l����w4��f����԰c���y־^������������}nw��ِ�OjB:�uحr�ܳ3{�����z\���G6\��S⬮��]�c�[DXZ�~��u�̙�����ݾ�,��_���5w`�am+"hwe��޿[��}j�?\&DF�/���������k�?��=��c�������ET�O����f�/N\����=�
 ��^����U ;u�T�A �("��AUN�W\���>��w���>P	�<��Þ���'���|��O�����G���G����/v��ڼ��s���]���_=�w����_�U@?�������**�~HTU@$��I���?����O~;�����������������?$QU ������������w'�����'�/��?W�<�n�v���Ǉ��?Ǳ�=��n@�|~˂�H�*�ʒ(� ��!
B @��ʒ$ )"H#
J*B�"H
H+"J
H
H#
H#"B�
@�"B�*B�"H�
B"@
B�@�� ��Ȓ)
H��"���H��
H����B�,)$�
@$���
B$�
B$*@�$�)+"@����
B�$�"Ȓ�� Ȓ�)*B��� J���"B��� B�)($	B���*�
B���B�!"J$)*���B��"B)*�$�ʒ H��
@"@
B
H	
H�	 $)"�)$)�)*$��) �� ���
D��FD��F ��\*0�"�$�����
��(0���

@+J�B�*�� � 
J�"@�J��$�0�(�$
����
2$�0� 2$������0���$�����$�� 2$�� $*���� $�#"H�) �� �"B$)�
���"B$) 2$B��B�"B���(��(�"J)"Ȓ�),)"Ȓ$)+"B2��
JȒ�) H��
@��)"H�)(B��)"H�)(H���#"J��	
H�$�� Ȓ$) H�
H��
B$)
s
dHF�!H�!H� IRV�$HR�$HBT��%aHD�!IRF��$RR��$aI	��$eI	��$� !HaI	HR��&�D��! I�$!I!HdH!H$H	RY�� !I%I$H!IdIRR�D���!%HdIR$HaIIRYXR$I!H!J�D��D�RdI!I	HR I�$�"D�RBD�� � �%�"�RHRdH!HdI%IHRdI�!�"T���D���	��$�"�D�T�D���D�RdH%!H� �&��aIHR�(R	!J��aI�$%H�șaH$J�R!H�&�R��R�$�"D��D��&�HaI�&�RI�(R �&D�RIeH�"�IR	R$H�&D�@&D�R�
D��H�"�� �R�FD� $a`aaaHXEFAFRAF�Q�!eA�Q�	Q�Q�	T�Q�HEE�Q��Q�XE�Q�BF H$a�Q�AFH@de�Q�AF dd�Q�RTFEXEdd$aA�d@!IUdHQ	RAD�@�$$IRBT��!%Mu3�@���������~��=�ET������k����_���h�=�:�~���~�������o�?���}�$QU ����~�������>}��������t��I��{O��u���v=袪���}'�]}��]�׸/������AU@=Ȣ����������������������`�!�ǧ�:��
�l�8}��@t��o���}b!�����ٳ���#F�~�@�v}�A�:EP����G��z��袪�w���9���y�i�=<��|����ϫ��}=�ǐߟ� �(��s��x?����������������|����t�<o`y������A�q����>ݾ�c��>8zw�z�� ����^��?.Ǵ���>��W��Ϸ��"��GLv�o�$=�I翼�w���s����v�v=���|����QU ��9��g��~�����>_w�QU ��y�/����Ӟӿ��������?����z��<���PVI��X*����6` ?�����v�� 4      P                  
   
       (   ��*��D�DT�(�"
		
JQ% �J$�$)($U EJUQUH@�QD��H��H�   zu<B@UD�EP����8�Q��xYE�p}�a���)��ǈ�p�� �N���U�wU��ܯ�n]W��y�Y��R���Է\��=��h  5E���P|�  p w0  ��"	\ �l��

p@4@ ������u*(A� ��{��#O�a�x>�|Ϫm  h �T
@PH� �>�T��t8���u�ݻ����n����_g|�vҽ>�E�i�����u�_;+�����@����7ҵO��P�]��緯�����:ؠ ��7ϭ�*����]�J��x$U.��ӛ�x��[���ˡ�:�����N�|�*�)��Z����R������^��}�y�U�Y   Ġ


�*���
���JH%�굻����=���_K�W�{��W�{�	�v�U�g���W�;��k��;�^��zg��@����q��uU{� h   ����W���7�R�� �Z������޻�L.�:�{������HR��-F׶��\����X_m�wN�@�(  ��R
 
@�P�RE.�s���]Y����k绫ke��Quz�����U{�ꕭ�Z��������ZV�wYUnwui  (OmuUWv�mUK��J�U޵��g�����������^wO[�T�IJ�wUC� ���c�`��`  ( ��Q��I�T�f}�{����q���U*p��<�l=�>�{�����pe�|z�|��
  >v���ב��;���r�P�ǟb�z�����y�w�h7��p�� �>��GxǾa�}    5?P)�*UM4�&���j��A�d �S�j��ԥT�M `�"~%JJx�  OT�#h�@� I���R��$��i�������v�_��<�3v��z����� HB r�:��B�� ��$! ?�!��� ��?��o����ns���p�\���w��qҖw��^�>��J��9o1��_���{D�-=��ޢNw�g�R&B9�����i��(��;��&�Y��<�m8��O�r{s�}�qy�9Y�j�+z�#7�3Hs�����-�t�`�_*�zT�F�/�	���!~0������{ؖ��zz�s4C6�j�#���������P�B��:$�E�8'�7"7ط�^}���{���e�N�����A(�����{n�ɋ�U�k�����#��s�aϵ�nw�=��.n�y�3��G9]�ܔ�-���97���U��1oo���˃48=�P%����1��C�^�S�U��T�Q��^�w�y�{�ù�%ޚ�B��v����՘g	0�醊׾L�}N:{bԻz�SF�+��ogt/Qpj�u]�w������]},s�W���x�=w���l�\�#!�:�4��}�$�2nQ��2�V��ܿY��c��l�� �sX��y_�ž�K��Ǟ�g���#�<�޽�M;y�ܞߐɭ4h�t:<����<Z�BJN�Q�û����~�8�h��P�o��r���7�n���}�ǥ��'�z��绞�'���B�����5]��Y���ŎPN�VO�[w�}1j[zvlSfC,�{>��[�Eh�c�,�r.g���=�G�[���R����h���Ǉ�m=�qP�b����=�|��ݾ�������׷��}ފ�>l��<�{(�i[�ȷ�.��g�{ׅ����a)@�c89�e/-)<�~r��W%���3U���S�Zxx��>�H��M�:�UJù���;h�y{�x��_a��Ʃ��}�W��{��q��6ZZ�s�G"pnR2�=����棭�B����y�����L��ݻ��!=	,R��hu�t{m�=}�{�{7���c�x�O�oǅ)�wdj�.Ǿ�r���{=���<�w/x���w�U6,��MX��*�9��5���熤��|��c7P򫜍bS���8xe���U�3��|�����vz��ú5�+j����������ݱFtݰҶ��g�����_0{3ð��v{Vw��'��ë�yo{m�r#ٝ��Ĳ�Z�J����;�ޙ}��2/�����v^K���o?Kf:������ם��걜w����K���A��М=�y{�Gr�]0O?ud�>#���P�<��7���)��Q�"h��{���������{��ۯww����vه�e�uEp{B���l����o)qq�{k�{�]Д�:{��=<Rf�O���y�ɺ�ީz�����z���|��� �'��'����M��>���)�⚟�����6l�����q��D��]��Jk�����=z�����{Z��B�}�j��~q���b=������f#]��E��yq|}릝��8�|࿣t;��}�$�;��^8��w�[<؋���_����t��Z����.�y��\�;�w=�g������n��G���: �ɽ|��f��}����t]��>S���nL��CWo��f�x^ў������R�jɹM��]���m�<V�y��U�齙���_���=��s^���s��}}�|�5�FM�]�٥�1��̻���$�ӟ��x��E3��{w�}Wn�/f�'Nq[d�=ٖ8wc��2'g�m�^T�����S��8�_�85��-ܯnU���x0��
�8&n���1ӗ���}���=�;Ff����D�F��B�|y�S}0ݷ���o�.���_9�w>:�y���xs�ńy%���t�ye�x?M�)oWa=�����wp{zb���7N���Õ�����1���㫵�����X�d������w�{k�T��ќ���*�n���<�G��`�:+w_{��Q�����}�"�pE/N/s}�猻�qK��#;��P������n�q�~�\g�>�m9�5��1��|���T}"cVf���p6f���}=������p{O�LVx�i�+Ο,���/�+6�t�ʹ�:0_� �s���p����:��z��q+���M��Ăq����ǂ���5u�-ƍ�>�i�u[�v�yk=��3t<f'q�!?�'8��op\<�-��w��#���Ym��}�{�3�.I=�h�ހ��&����}����>3�V�7����(U��/S��.ÞSY�-���ԽsȑPѓ��(���m���{71)v����9��ϒ�=(����r{o[��e{���o���(�pc����=f���P2,���������K�����k��V�;���e����y��_z��E�����i�������N��;"e�QOoT^�ٔࣽ�3��i�f!�z��#��J�K���g��q��M���F~������Şx*��t>�S9����c�W���G7���-_�B��)���q�}3�\��������2�wy�^b�ofoh~ѾthG�~7P�gm�8.�f,�W�9ܳ���{�2o��>;�����V���'���ٚ+:ڰ�_q=�M��ض��;���L|�]�9'_n�^/g�<���q�OY�^O=�=�=ᳫփX�w�<��uG�T'��yf�py�W�XO��N=��f,�1{v�G4�����|g<��yz��Ǚݎ�L��ﻷy�eO&��מ7^.^U�|��3���ٍ�g��/���=���a�t�J^|V`�v�5s��t���'��˝�r�^v��K$/�j�c��	�T63�yy��w��ڶ¦og����l��=��c�w���e����Ky���ڞ��/���n�hOvzY�5�7��9w���d�Ҝ���.A�N���ELW���Ҹx��JH��K{]�ӯ}�||/��}铜#ٙ�G��nM񽹼�x-�ﳳi����������?u틓��x�y��-z��p��^2�47R.��ۓ|}��5��j;Ĳ�#&Q�;����,�n��xq��?oT�l�yt�ͬ��w�n:�(]���e�RS��Ey�%��۫5�i���b�;�=�r���ܶrџp�C̝�"��ٻ��C�<�x�^�+e�mm�Fn][�}zzӶ���_��fS�?!��q�����j;xIɽ]K���;�d��n�k�3��D�7%Qyy$�mLx���1�;���<��HH�'3�4�<������w�����|�m]����x�P�[���B%;�>�G6�фgn��0?N����gr���E<��obpzw��9�v��Eeo�v�O�L������oS˲��3Ϗ|\y�)��x�bZH/;�蹃�F��m ����ŝy�h� �s{��⯫^I�N7�,��y`���T��rNҝ�AIy�����oۛ�+����&ў���f��ڽ�0v9��k��<�F�^�罼$�q������9���o�.!1g�����wY\��]y�o�{�Bu�ӌa�Ѵ?o��{q{����3<�b�_j�-'p��s�V�v݃g�ދ��`ˮ��%��w�5����z��ܪY��,c�f�kfн���o�`�Ni�����Z�Z����o��d�����o)�4LÛ(^�zYw����ʳ��9x��n{��7��u��y���ٽ(��s�Z�{�)���4�m۝\zʼ&�p:D���|��f0|���x�����������w���	���{ۜ搐�w�w�r�0�{�D���_C�s�}b����9��]��=�͚X��M~��?y�W}ٓ���\y\�-��{����ے�|�x������A^��W�����)y��T��9tz�w��w u����WE}���7�������t�l��C/���h0���z��Ӱ.������ۯ0�g����k���z�U����jc
��I^9���.��0d�m͞�w��j�Q�x��{��r�k��B6���{W_m��q�[��W6]�vbݔ�Ź�|�YO�c}4��({&7��^C�7�Z���V�y�Z�D
�s-�j�ٵ�J]Or��Ϸ�F��)���sOh�I��l#04��t���5W3�^9sӽ|֍���d�W-�]��M��@��#/�����8ٹ#����q7�	ls���B�����f���6���x��,���"���~��G;N��v��Vu�����k'#E���y�8������ǣS���뗷�F��vܦ��|w�_k/(]�=�n��G��Z*rZ�;�99��d>�J��z��J>^#���Ǽ���;lx�k���A�>9�)9��>�|�|�,=�߻��o���nY8!�_7��z��e:N��6[|��ۓ{=风��Fc���΄=���	����Q�[蝥�빞�g��$(�xHU��z�F��������!��{^E�x�n6�ʻۦ���{���3�`��{���K�׏r5���:a�#x����ar�E ���6����>���w����15����?k�9�����{ݚ������I�"���6�t��<b@�Y�}&z�_�PS�������]�ܚy�yq~�L#>�PFo����>��S���t�ᕑ|�Eݻ�.�yot�5k���E�}�}42�G{�G�{`R�Y�{j��lQ�b�=���$»7'��M4�f[�p���(բ�ͷ��O����7���rɅ�������5}��y{t���9���	=��ݭkŵ��큍�<�t����g��h�K�^g�΄��ε�[�G?j���Ōe�<�n�\�����n!�/-�	7�����V�9}���ݹٯ-|�D�:/�m����4{��E����ِ5���6�/��(Xd�5�Q�Ź�4����/3e�E{�-6���}�~^�A�n�O{�W�43�5�^0�t�H��t&y	���/g+�g���زe}�s�})bG�Z��q��O!��r٫/p#�s��-�6X=�7�47|�D�?,\����}�xg-a%��uz�sG����v��s\G��!t�9!�~��`����C1F绽F}Y̿?)�/��~��"��k�(���opY���+�=�C�Z}ϳ|o>�2��N-�{ͱ�ʰ��n�����K�̹�?{8j�Bt��s�m��%>�����B��8��h�0������rq��+l�!�*���{c~��O����f�i��.q�+Z�?����,fu���sg���%�V�����N��鏇5�3��ڤ��O����F)�����W����{��N�zӆ�f��uu�\+�pzg����uo|�]��<;"]����V�l��:��8?�5�3����ǓA壙��z.��_�x�B9��C�>ٹ駞mu��=�J�\�H��m��4rњ:Ai�|�����z��-t[e�M,��Z/�8��3'������F��sw0���iÏ�8�7�ݳ�uZ�,���H���
�[SB�'���p�K�;��7үE|��Im���oplQ��LK���'��_���M=�}��韃(>ߌ�Y{[�&^���T�����s��h:=Ҟ��3uu��{�w%��3��m��y���K#�����z�'�x/5�fI�=���3c��Ϗ�o��W�}W�yX���Hկ�&we�I���uS��`��\�B�!�d�3��sƛ��:{���Ebk˓�̹>�7w�'cE������j��qe��)g�{><3�輟+7�{�b�ءߎ���m�g�{})Ul8�JG�:
�۬pu�o��fU��畮W�a������x����u�Z�ٺe�Ӄ@�-[wg���xG=�6�q����`�Vr���<���j}�>U9'�r�^��f��g�z2۷��������aP���{{�����3�f��އ8��ZVsì%{�;�Y��u��|vw�3����ooo=5���1.Y%����@�|�g������!7���W�M����38OAQ��0T���X�����g���G��r�A�w{ٛ���j���ǽ{s�wir���A����^�V|�ٯ۽;���F�I�7r��r���;{��L4��H�@�r��z|'rs��	�}���#z'�ȅd�����Ƕy�ٲ̈́7�7�wT^V��ǝ�9�z�ק�T��T��١.}=�Wd���A=���٧xs��z	�f��T���E�=�_h�UAUw����/&OL���}��� 7N���e���`ln�:B�i^��qv;�Q��oa�9�����*z=����N��W���白2�Lv�GZ�8�H��֝5�=���8/�׻uͼ�CXۀ�P�Ad��}fb��]1v��v�7{7<�����F��=G�yz|�q-�f�VF\���p�]���*���]*ɽyя}٢A����.�����8�b�p��M0�Ȱ�g�K��,1�<�͋z�:���0)��J����BA�^�6�9k���=���z���[{�էV�����?L�Մ���Uǚ.g<�3ٹk�I�}��n*W���'�6l�F���|�}��|�9��zr��=����&�]���e�b���c�r9G��m���gn�B�=�9�7��{��{Rf��F�y޽��ˈ\}�\~�r��==P�_f��vn����=�����s	L�'��~J��l/nE۽Oownbל���\��<�%�j��H�g���h��=�v���٭�����7ǆ-%Gٜ��F/��I{�<x�H`�!#�76�C�l�_d�<q�By7�v�q̽<���On4���ĵ��Z��������{|.-��{T�\g�~�^����7}�#�Ch7ήi1}��<�y���yFv!��琛��ōMwX=[V:��Z�sE�o�v����4��F��|��������͕f/fi�`�1��^�<�����R�l�y�9��zٕg�Wi:��5Fz���%R]_����c�Ov0�^��Da�o��4'�.o�zB|=��FO���[~2���׽�Hv{�Kُ��{c�{�/z���h�k�X|w�ݣ	��X;�܊ͨ!��%o�]��cŎYl�5z�x�¶z����zul��ͻԑ�ZP�~�e�trǌt��ڙ�͞��-cr����M}�{ƾ�>���g�3�y����{�_m���i�aS�}�ym��?/F��Ιә��;�@�z��(��Dm��O2�잯ܰ{��ٱv^�q�pǞ�چ�y	]�j��1��٪��b�����=�a�Q!�����N���bǬ�=s�	�}���e�"����%���z�)Ny�J7�����r�n	�O��1y�Ԭ��W������͞���7LQ_v)�`�t/ �Ιq(}C���p!����g{s1c�c���4�n��n�����g�>����w��l�9L�>Hs���}&����SrQ��3������X�v���b��7=�s�x�c������GU�b�?cWˮvY{��{�d�IUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU_�|UUUUUUUUUUUUUUUUUUUU�-N�$0�Ԝt�l����{���|}鹾�LvUx��Gc��YK�wh-���cvSۅͫ�Cs�q����-͏� XK3b�.�5�[\dY�J���ԁ�A�l��A�-���g5c������3������|�y����n�-�F1���U���MH�;0w.rPL$0@h�ںU�d�/]+�]ٟt75m��ƙaqEGgC��!-�ۍ#"�F;2��8^����.(�1�nk�tM[�cG2�eۥI��r͵���ǡ�l�6�t�(��q4��gO�����W��k������^��+,V�rn��5�N�e��W���*[��;�b}�[���sv:�H�p���/l���wax%��gJm��<P�5�k�]��/�m��iK��l4�&.�eH:U��M��egyd�Wq�nɬs����
�^@�7F6�t�O��)F�z��v�z�vwK��\�<Y�Q��Z�/��K/l��[�T9�eKq�o.����s�	)�0$p�մ���y�Bhq��k�Vʗ�ۮՅ��j7V�;ڪ-�T���9����jM)�闯m�O[���h��4�McrG�����5aɲ�6IB��%X���:i}9��<��w�)�B�Ml�,�T�Q5�T�O]���ڦ@��2���K˹��Z�vkv�!mt��U@���L��[��F2^a^��)y"��<�8��i}d�[�w4���ƻ/����i��9� e�����*�Q4�˶+�"��%m��WX��+q�Nh�tf�� �(B�;h-��,������vt>C��ۋU]�dt���	���<f�s�w\n`�&�r޻u��<����r�2�5q��xzī�ۉ��\�Y7B�5��Y��������v6�ŶN�(n�Y'�z�3nm�=n�Z�NݞJ3�ջl:�kc�vW��4�h�q\a���p� �:�b@�*-ر��ͫ�qj��l�e���
��/1Ct4������tk�=L[<f;٢�¢�߇}�E��x�J7i���p�δC���v������L�n�p��K�T�t���r2�9�4Ί�Da�p�q�.Ud+t볛�*c�Xwh��ȡ�M��رcj-L�''Uճtr\Cvl[��q;���ۥs��h&��R�Ʃq�gn!|ufT.�=9��k�èh̎�0ѡ3�q�6^ے�n̝$�W.�m<PY�jz���i���f6���Y݃��m�nu ͳnni�ڕ!�l�f)S�fv��p��Dˆe5e��+���L��	�I�m��r�g���wQ�ʶy��vC�<��o]����H�i9G]KmNp=ԩ�sJi���]�i�l�ƞ�i������ˉ�Ͷy�G��s3K&�E�Yn���p��^7;u�mI�U�������1��*��p]4���+Ҡ>�\��&B���v���'nuه���g��0B�Q�uOan��"ۜ�c�L6�R�:��	a2rƶ�(�ant���9qlQ���Q��)L���$����qo��;/~�0/p���w%��tSFe��4�mr8f)1��:Ύ��rkf^J
�iؗ��u��y�W>����=cs��'g�\u��L��%8�b�v��Ȗ�S��..�A=b���n�{�#�������������mЫZ���	�Se�X�˒1ˑm�kx.�X�8l݆�ͷ@X닮��Q%��F�o׋�r%8�18�Cr�<ou�����u�� ��i��|g=����6��{����5qm�bd����01�/E�Mt����X�-��W���c��k.��	�[��B�X&�y�f�YatuQ����k��%P��㞷2X��v�g�n�cX�eY�-�+�3+X�2��A�yl)����7 �1��� ��M����V��ٰV�R:
L[efx��,�u#��T�SZ�Ύ�fƅ��Ez����>��M�[�J�g�3���l88��L������5�.�n�QZƓ�gn	}���k-�<v���Z2�ea�`�dHA��c�nunڍ�
�U<Ɛ���]�<T�u���3�;7��h��e��1.Ӟ�8^�چ՗kaf�$ct�s�,\
ʅ��R4YI����M�`.M��z�c�>���pqݱ�Y�G��k��`���nՃut�PУIt�+s�;Kq��l��Rˎ�	��m�@��s��vQ�٥��7<��@:��G��{�6��6����c�rp������Z{Lm��l/g��X9:]�������>ˮr���	b7VぃE"[#v�z�\\��a!X��k4�Zj���P�9��y�h;>c���u�:��G��:݂V��ȕ���ۜ���vPlfű�[>��c+'g479Ẍ�ቇ�X�&
�zm�qn��f������u�pN��<��c{<�TG����qZ$�0i.�]�lDsۺ��G��{sv�X&��w�q����xr��p���f�v�Vx)6N�Ϩ�ٶ*Y�v#ug4�Қ8r�m��l���r�5�i'"ܛ8��7j[3u.l!8�@�.�׏�����lB�ݷA�O���g9��ؽl�el��<�bF!3Qx[�l63l5�e��h5͒�L�+(��)d�P[���{���}�\� �̿C5��ӏ�1-ۯ��}�C���X�	��E�v��̯C8�;q,[\u3�t���im׏[��1�3�ܘ�ݝ�6��/1b����EjVw�\ݜ�V�N۸����ԡ�w3���t#t��CG�+�f��Y�K6�5t�VV2��.7�J��(��]��j'���.d�"�mm�o>��=�֜v��k�e:�]�R���4q0�Z8��ݹ�F㗎�����KZ��y�������u��˫���2'�=g�ඳ��Zѧ����]��l$�A6:��d�=g��=������۱ι�7�����*H]�K���e�U���l��(9\�يRE�=8��u�\�gnږ�fkp�\iV�5�Ķf&��-�֧+�&i���4ҙ��S��E�VoV�OKn5Y��n�C<���㋀3�.5rjRa�KXj�t=�Ӯ��y]�p;G&4��i�w��M��̦ 6r%����l/�uȗ��)�x��I���w�E�g4�3��]_��-]����0VQ+jY�����p�5Qֳ#��-X��lݒv�!=n8w)�Y�|ú��d���p�]OWWm('�<�0�.ģ��V�a��-�-qر��;�f��q�OA��kmbK�STWg39ݍ�1�=�HF��$JpCk!�yHѴm'76ތ{p��]q��T:����`�	Y�5w6&�ӑ�9Ӄs��y^�,�3�X2�u�#\e�c��v.3�pn76:NuN�X��x.y�8�=Ӟ8�WZ3�f���ݯ�>NQ%N���������Vx�mՎb�����G!���У���;���vDC�s��.M�N��aㇱ9��)�sz�K��ulTV�Jv�v6���\�%Ϋ��˞�Oi�p��c�mv�� L��M�՘�F��5�vX�M�h�t]U6,P��H��[Bյ��sj���uK�$�k�0�U�fmIn�."ڼ��tّA���q�u��:K���yݣ��c�����˺�c-5Y�b_<_<�#P��YMn���m�Z���ax�1Z<��ո���@C88a
�h��͚bfh���n�D�1�76\��7ђ�erqX���4�ka��p�m=���+;pyz��`�k�l�*�i퍛����O�pn^�mcp\�gl^.���P_6-u��f�(�s�7���ɛ�w�{oKF{2��v��m��ҰWA�m ��s�Ё����t��5qi(��Ћ�`M#�>�]k��r'�Y��Gq����Fi�S�+aP$%t�F�2�g���)�r��4T�A�e��s/N��N�V�m�뜝M8-M�p:I��އ�y��9�7[�n�>�R��(�&v�VŪ�JX��k�@,@��\��MR6����6q���n*7�lfG�� Υ�2�=�v�>7!��y�l�.�;�K�ֶ\:����	d����|�r��n�f���:�S1�Ps�X���ي�}���s3#���yY�i��&ME��+u%��!�V�Z����/����[J�1��pC���q�ݭ�A\���ӏ6]��빓Bڵ=�ʈԆS���r�=q�4�`�;	َ9f���*�h��θD��m�]��4���M��<��Gl�r��:���:ۛ���ʹ=k��pLy����Ip6Y[]�նSE��]pk��du����Ĳ�M�,
��-�M1)^STr�k�j��'��,�m��Y1j�kp�GQ�����s� ;��n�uuw�ɞ���Oa:뭗�/��n�Y
�z�wJ��NX�㴹�5s�}v{�b�Q�V#65��<��֊���]�$ܖ���8Ԗo;iD�U�3F᩶t[
T�Sղ��g�q6�9�u��5�0��l�tq���\d��D��5<ժS2d^C�5B�v{����:x�)z�fۡ�u�񳼋�����瘹G�oN�قX�����"�+aV.瓇��>t�䧘BfkYL�wh+�o1�v��3��ٷl�����ܕ��3�.�,`T����.�����),�5*�W3��2���A�t����:�ӣ����囖̺�F1���l�3	�5��Ƅ���`t�� ���t�O���n.f���؞:=t���c�4)U�u�.�+iZ3����K�ؑi�.���i��o/��Ҩ�-�o[�z�Ds��YX����h��%,\s[���;�9���V�fo���6C�}�FH�^U��;��U[��Q��nN5��X�ǀ���v��Zs���Q�\�;��\Zs�-��mu�A�'og�K�cr�/L���7Z&����R�,9�֧�˼�lsKt�Em�[ji!qݟ/'�ш����Kn>�Ȥ�hUj��ک��l�Զ���XXf!R-X�b�qV���
�S��m�����$4�sӥe��<`�����af�D%_hn(�[ugs�box���6�.l��XC3<�ذ�1�'ogu���MLk�x�kL��b���^cG���������4�6dneqlJ�Hn�׭���oGn���^5`p�Ans��qw8g� r�8�8`{"�ue�Yq��E&�MkE�CK,e4�,jkt�UJ���\Vnۧ�x�.A�ۥP<���n�����]�<H��ԧ68�OM�W�/i��<p"�1�� ��8��q��@�<:{���pղ�p덴�u�l�]�fkL��r2�����9$�rN�@�I�I�$�O��������5��#�_�i�{�kT�_ɬ"dq��G���S�k�+э/�%W�L,!�����!0�����d���ΐgڎ(_/9��a�)G��&E�.�bx������?j�~�^r�F=w�n��"���|<۰7�0=�a��yJW��!Kw�xb�������Q4�9��u䯵��4�iӦS���}��9�P�T����N���g�sL��f,�^>��F��.��t���p&B�oN�,D����ꟾY���Ba'���{7	��A�����ʾ�y���fI���ؑ�-�]�6�%�r^F`\q-y�>�J{|zy��#�n�שj��[=v1�*�B�LC�"#Z��ϜH3�<�����pJ�ˎ���kǹ�y��!���e���BA���=��<���v��#O{�:V��dX�c^��k2T�a���ᘵ8���;1�i��[�#�l���׎{ݏS�D�>$>xr"p^�ο�m�jH�Y�؋eg���al��O{2l�FG��ﯧǸ��;KŲ<��[������y�m_w���iK�;��7fF]-����w3�vw�r��ܙsEҰ[�w�Լߞ�h���j���L��E�bgq�R��,��>������'�0K���z�Fo/{����ȵ_Z����.V���t�n�I�0������g�Ʈ����	:�$n�|�-C�{%ϸz3���^����m��g�ygi|�/Gqm"B�h@�M�N�>ƹ�I$������l�����5��S0p�[WYb	�,�,�:�m��J�l�M��=���
!����u���>�D���yE4G����ԛ����n��r8&هݻE�f&�{2g;4x��9�nԚ���-Ґ�9[��:g:��v�1�N�-�U��X[Ŗ�]Fm�p׉m�i�T*���i�h9��bX8�ಮ7��F��.���nD6;,.�;��
݇�7;<;P笝�x�2$�^�n���;7k��/��r�#�kN�1�*���ǆt6h9���
Ue��Tt���5ҫ����ָnl�Z���uW�:�hWn{hB���Z넸]q��n�I��������(���c�:۔�,��ulz�Wg��v�ǜ6zؗe*�{.�.�r�{��3�8��r��N�u�W�n��5̖͢�8WB8�Zi��MZkv|{��c��Z.�Lˁ�:hJ�zf���^{x4 �����J�`ڦ"�K��a6t�`8F�d֔5e�]�T�]lq4���2�$#)�W�+�m��rNF�h��q�>��Я:���R��'n2��*���6�Ch��6n�� ����W����3ާ�ݞt)e�.P�m�W]Wݮ��k@�Ln3</<C���X�ckR:�n�dW30\�-,��(�s`�V�t�t�6�G�m͹O���8�lr�UV+u�[؃��u������$n�Lh3[k������y1�<����:���k;�p��fa�v���93U�a..j�F���wM�����N5�ڎ��8�M�7E#����)�H�+�PMt�6���q�͹^3�p���	�1��K&��!���nZ��t��t�.�l5�U`�j�k0]F�0��f�Y���>3��y��J�1�10�e%�MmR���&��F�벚��NU�'Z�۩�c��[Ih�e��bYt��U�fa!h�n�6�Uc�ns�.�6l�Ti����;����8PUѶۆ�a�A�ị��Xk��.%�[m��X�	RB6X�v(q��E�&��C/�q�B�	���3N�,$'��GKaD*�ms�Zѫ���T�m�9��0����e�eí�ӵ� G��S@F�wh�X#[�LD���j�4�;�IG�}v������H]M�nv���خ1��O���Ϋ�,=�qC	�O�X��GU��Û:��Wdu�v��]��ٝ+�Z��vv��]�.�cj�u����)ս*�0n��t�y�6!���K��p�545K���y����wn6A���u0���M������Y�=���C�vՙ�Lkԯ\���p0�։l�C�k�g �i�c��s�����#$��\]z}(R�ȅԣp��f8�9�.:㞞��^$��S	��YLqas�a�^�C��9�#}�$8��)z��3�.��Q���1�-H�0�?[�Z��y�T-=�d/�1ͳ/�$�	�(q�]U�x��2�	I$C)~�j��p��+�g�چ��8�8�׭�:���?a�}��-�	��(S�3!k/�$b�Kw+I�Za��j�4�u{p��%"P
U�[���	Ȇ}�i�s|p�?z>�:��O�ԅ?q�����Y�xΎ�� ��u>ڕ�<"���vƶ�m���]Yc2��	n��c�1�6��JQ�U&�2��UL6w�e�Y����F�-ys^��4ڳ#�q��OU0��N}
P�\,�O���xxD �$���E����-3JM�S�Ece"wtB���ӗK3x��KO���?��ك������{���a�O�f�I"D�N$�0���~ϑ�)�4�8��-��c>yuKOiy
���G��q�yN�G�]�3���P�F������㇎�m�<��ap�#Q}Q��a)������YjiӕVJ���˅��[,b���S&�ic�'v���rV&�����In��:�`�4e����&����g=KY3(X�[*H��}q�Ч#�7+ϰڇ��ʥ,�?U�NZ�tё�.X�4�*&�?q���_,�#�E�}�48᯽~�D?B�]	0�� b�C���i�}��4ڹ�����Ϯ�y9����2,?4�҉5ݮ�.r�w&�Hh��X���0*9F�����#mU"+<��n�����wU�YN�Fp��5I$	��C��qӞ�NR0��^����)֡�#�*�XT�8�˪ߑ�|��L�uCM>"�ゟ����)�Ec���K�ZY�k�VŇ��ձ��g�ڵ�wQ�R7]��V^�!��ˇ(gA��R�pg��Vh�v�.��l�2j�B��0Nݸ�@�,&u�i"���MYji�q-������irI�#�'qe0�0����"p�����TkL�L��a~�\,%�JkP2Rl��MĜ�q�8��eji�*�����'u��p�<B��[C���v�m՚�%���I�'�{�4��L|��³\]̲Ţ<��ƀ(�����k�Pi"nrRb�L�(� I��\h��^�.�"@ ��"���Z��t�`[�&a�\a��0q�����yK4�ըqm:q�U��~�e��0���w�7�uN�1f�����3��Uv�FH���˺��ny��������9-ӎ�)0Hۑ�ߐ���*a~����t�wT~�1vmyN�F������i�2N/��C��l��i�	�˂(���`�]��O�����N3j ˑ�T0�ƽs�-=��-c��Xło.��p���)~���()2bb�Q�X��0OZ�"�Cp��vPib���ɽha�Lu�C��w�|����Ɗi)R�#L#�1K�q���Ӕ�?`�ۉ��`��m_�nŇ� i����I! A|��8��k���w\���E��(�S3]��}��+�\�( B�I{�|Ut�v��4��=4Έ��A��*P^��@�ݲ��'Zs�j{s�.�.�rA8r�9����z�3����s�k=�f�l͉�[-�����FX�0�_m���z}�V']��z�G+��������N����[���'��9"wJ�uɑ��0����]����-�w9-+�:Ʋ�����@��d��D>�77��vW��3՞�ฺ"��E�ڤl˅�j[�䕬�.ыZ����kU�]d���u���7�񣷷hm�zX��u����8�d�/�oO`�\/�`�#.%i�/!n۟��M#���C���y�4"������Hg�/�a	0��9�t��چ�kXU0�?[f��4阌�$���d�"rB8��5뾙N�F�Y�.aif�ܲج�V�",�
�ME�^$H��#ϰچ���8�л^Z�4��b����gY�D�=��[<Z[�Z¶��,��~qlVzǱo�)�i��V9�A����7Ǆ��oݧ��L���u�.�5�Y
��T��4Uԛ�Dh���n,���%Y���U��k]��g���O�W�
~�5	���0�<Q�i\C�oeC)~��
���n} EH��Y�m۫� H� P
�ÒN��ݑ4�ԁb��C8c��,k����H��"`ez\%���mC���.0�?r3�Ψa��W�L��b\���B��"�*9��/�&ܭ"�if���ج����$��G�~ϙꇏƐm���5mI����m՝P�N�srAO�s!n�:�`Ńu��.�ici��b�.|cI�FR4��ӬI
p��%���p��ei"�Ӻ���ibe���.!Z� �r]��V	�=�ִ�^< \7�L퇶·�ֹ�g<
7Y16�Ƈ���9Ӕ�H��1���:����P�-�%2�0U�6�,%!p��T4���)�8��շ�UӠL����u�6��4)Ј)GL2���G��]'<�g޾���)z�R(beEݺS|��W(�2I�.[�Dsr�H" Dl�@!s�(���d׷q�k,b
�M]%����m��t�R�L#��V���eȁ�Iϳ�/�`�х-=�\-��ql���GY)�p����e�Q�$G���%	�[�!L<t�Ⱥ����x��R����][p�g�3.�i�3!O��UH�Sg�Rٌ���-.a�Ea��{<h�l��xͻ�oQW7N�v�ڭ�1X�VG������k�Y�$��1L<t�e�>F�<m��ڑ�Ks��.G8�8���:���2�xЧ�7�������+��i7L���%T�ƪ�ΓÉӾtO�I�����cp�ҝ�t�i�u��/�h�g����증9��c����t���Cs�Ҫ�k{8[�B�!��A�h�����3���7���ĳ`�IPdLB�R "#;��݆wv�"f	cFnX��#�_4�,h���M�c�>��z��ӄq��9j��+9�?q��v���x�.��hX@m��k�h�'6��&᛫��l�$��wGmm"�r�;����}�7�v� ��yr��٪0��űQ�5�:���4�V�/��CƵ^���GZM:�	Ɣ�[q�T4��XH���:vٔ�i��R)X�9��a�Ht.N��N��n�<t�e�ϙ�n\֖-=�taz�|3w1�-=��'[л���E�j�վtN�w�>*�if��*ذ�m����0_7B���C
�V
C-�DƓn8�~�;�:��N��kb���!%��,�}���?=~;�|_c$�X4>ۥILĖ&i4b��$r�7wA�#���6$��-�\Į����Ɉ������}}*��S:�ֹ�9^1�is��1J&���W9k]�`X�l�]��<�Wy7�!�Y���<���v&
�97h|D�Uh�n�{q���c���H�9��y���:$\��nC��/l&�b��6�7:�$�������w���&��W���o2�k;&��X�1���j����BX��Y��c�5��0�CD��[X<�Yn�IT�a���̛G'3�&��a�cr�8ʺ*�k�Aٕ�(��k��k�15�����j�&ǃ`v��K��V�ѩEI!UP��Q�vUT-,��.���i}�#�޴MY�t�^�$nHʈ��Pq���;9mYK�6a�&M���z�*=����K�>=%�};����T[k\�q;�>'aأJ�nmͷ
�a��Z{K�=�h�t�<`�Q&�$`��qBe�-0�5�+b��O�-D-(�N�Y�6����G�#���HQ ሉ �9ji�s[��ӖՔ���]&]���~qlXz���%� �L�
\`�nH���4S<Ogf���^��r�c�G!��ѵk�BD�-
p��/M�g�چ6b����i��X���^��xF�P.ٙ��O��L}�>'�!FL��!c��gn�#��N}���H���0$�7��,���Q2wN���� c�E�d!4���+M�୊�X�媅��t��g�چ����W�TxD ���&{��
����;��%i�2�n��N�G�5u/ㆱ�_�a�D��-���i���)��H��Xϡ�+�G�\�-Bt�JX�a��j8L�7!��u��2�4������8����e#Oк�i�a�~����Y���ۗ�,�$ֱo�^ݑ�V�6�.��^���(*��.c�Jj�*�؉�ӎ(�ϙ���8�8�׺�z�X�*Zʁ3�e��/\�(b��#�A ��1�"��r!�O����a�>�x)���`�x�W����.�ӄq���5��@� j4LiÖ��O��B���BK�e,��|�_$�{�R�'WɏA0�X8[Aa*őJ"�+B�i� #V4s��ROx�����e4{�N|]��}VC��(S�(���O���a�[�`�T:ټtH��L��7�\�)�����^}�n8Ifb	�23��{��~)]!���k�Dy&8op���ם�����~�#���1��f�	�����q�X?A@�w�{����P���->T\�q��QFRg�O�z�zm�g<����u��0��>s 3�8>l4�����}����"�)8�d�G���sN�y�s�ac��y�Wl�r��t���h��T�b��[z	'���D@�ќs��}<��NV��O���f�<-�p�PaF����`_a¼�؀h�������3�?�x��C��<�A�LY��x�hn��;$8�-�4��|��<15�=����j�y�	�3�ǰj	�}�N~��c^�+2I�x��O��{Bѷ��3r�71�!��SEA5�������`)%�d�=�N[��D��6����_�a�n<.�f%��>d���7����{q�k�n�
j��M��m����z�in���k8� β��9=�$�R'�#�Y�zWڝ�Z��U[>��y�y��dĒx �'ߴY���h���烁��K�3�1��9���f a	�҇��L#|�Å�毫�^D}�}{�X\ ��@@0$h1u�����0Ł�D�&A1`2"�%��6��]A�]�dQb�bۄ��AM V�]y��*C|ֈ)���+&����He��`�Y8ʐ�oNj��r��r�I)���Ns��*C�H)�~�/ ����T��Z ������2c*C��S���d��.<�H{5�
q���ʐy�d�)�
�`�x�''��Ӑ#�~՚ԃօƹ��:�VO�Ri? V�w� �y�!��D�a� B�w��k�����@�'̩~�K�S+0��eH}i=���������h�� V�ߏ�c�ʺI�lSEV���n���1s�ǬX�:nrB�f9��e6��6*�2k��ӷ��'�R���@�'��f�:��ֈ)�a�+'�R}�u�S+���T��kD�{�� �@��������+g>��LeHs��<�Xu�d�q�_��n���+��������@�'̩�o5�p���I
Ì+'�RZAL�w/ ��ɦT�f�AO�+���<ʐ��`�Y7��ד�f�AB@�1�d�*C\^��7[5vo[�D�ֶ�S���d�*C�ֈ)�{���:�VN��2�
|�X9����R� ���+�VO���k����� V��T���0u�
y��
��T�֐S�L�3Z��7(�޶��X,�eH{5� N�V�\w2y�!�H)�
�`�o���'R�h�� V²y�!��^S9�Fߍ͚��J$aL�N0��s�I��6@ �!$0l��N뙜��T����I��_;sz1����Č�ڭ|��S�g�8Xc
ɶT�ZAO�+u9s��ѭ���R�[��d�T�9�S���+'��N�2�
|�R'̨�BC���Ld6�y����w|�8�{�'�'�o��~a8����#��.��㫤J���6��p�ڮm-0�>�3W7L�lj3Y�c0��Y6�SE�ev�8˓������AO�+�
���!������H,�eHw��=��<�1�d��!��S�a��w���T���S���+'s��'Ri6�R'̩{6��[iv]���l�[Mo��a��̩� ��˙xP!�L��h���+�3F��LeHn�
y�Os���u!��S�
�VO2�5s�]p���R@���T�;�S��.j��֝�M]o\�1�d��!��S�
�����&2�9�h��@�:²~���9:��H)�HHT���*C�5��
y��
��T�֐S;���:�Y6ʐ�ֈ$�$����)}=���V�·�Os̩ZAO2
�Y?f}�ru!��S�a�+'�T�}��m�<�R'�R�Z ��wپ�²q�!�� )�a�}�Cl�ʐ���
y��
ɬ}��i�in��ѳzַy:��H)�H,�eH~�s���
ba��̩���)�>�NԂ��T�f�AO�+s��<ʐ��H,���Ó�f�AO��0��eH'�Z%�`Fd����W@��~�n�̔	`�2B$�؂Y����ےi���O{���]��
fqyO�_�S��bm�[�^\X����d���
;!��@�Um#,�{X���w�k^�ŬXx��[>�S&qˇ���z�ڰ�m�%�<���]mxB���uV��c�]�K,���b�h��%x<v2ƓB�m�����v��2Z�16/ۇ�ݤ}aq5��K�&�&K��.���.٠A�ʈV�ڙ��k8�w?���S�7��쭭��]�:#1l������9�҅��Ͳև͚� �D,�0jVW�t��2�[��ݱ���I�.�L�&���`�R��N@�Ē�X,�ʐ���7����u�0��eHe��`�͜�Ɍ�oZ ��+����g�ru��e��`�Y8ʐ�=�wxAO VaY<ʐ��
~�t":��uJ�[xX,N��35�
|�Xfk��!�O2���AO V�=����C٭S�
�VO�R~�]w�
y�X,�eH}��AOuϳ\�1�d 6ʐ�H)����߱��f�/�l�r9Ӕ��5�
y���dϹ�9:��H)�
�`�u�!�}�uxAO VaR�eH}i9�eǀu��d�*C٭S�a���p�&2�9i<�X,L��p�;����W[�����HfkD��Xc�y� �y���
b`�Y<ʐ���?s�� �aY>eHe���|﹮Ad�T�w�S����
��ٟ''Ri:�X,O�I�w��~���@�$5Yo��'H�VO2�>�������`�Y8ʐ�ֈ)� %a��8��̩�AO V����HfkD����̩�s�S���d�*C��DI!�ɗ�4n�&�Å�����V6�r��{Y8
�[��"09L���u��혂5ĳ0�-Fe^�²m�!��S�
��g��O2�9�h��@�:²k��ד����@�'R���v�"��Xu�d�*C�H)���׀u��d�*C3Z �P+T�r�un�Z�{�7]]<�<ʐ��`�Y7�f^N�=��~b0X�K1�12A�~92M�n_�̂��$R
R��)�̄��F�{�d���1$1L�b��AO��0��eH}�_��S�`�Y<ʐ���9�}��a�+'YRi? V�}��Y1�	{ֈ)�
ì+'��|kZ�[u��vj��w�����@�'̩\�]��
Ì+'�RZAM{�f�X,N2�=��>@�35���&2�;i<�X,Of�_<�H{5�
u����T���O޹�]�,/\y9t�R��$
���h����k�²|ʐ�H)���̼�Ɍ�sZ ��+�VL����ԆZAN V���8�+�S��VO2�>������kvݦ��v��K�n��&�R�h���+�^��<ʐ��`�Y=��o��f�AN V²|ʐ�߻�����X,O2�>�Z ��߳|�1�d��!��S�
rNst7��:6l.��-� #m�k���g�3��\�m���kiM�d�l3B1pj� eRy��㔜����	�
������S����� V��T��k0o)��VO2�>�������@�`�q�!��S����o!�O2�;i<�N@�r��뿓76�mr�.w��!��S��0��eHg�޾o)䐕��d�*C�kD�v���u�0��eHe��a����'�R�AO V0���?f�:��H,$>@�'YR��ɭn������o' OĒ�����:r�>�����������f�AO�+�^��<ʐ�|"1�$$" �]2h�)����s�׷S4�A����$R�d�"���I��
bȕ�{��-�$4d�ؤb ���@�'�{�y:��ֈ)����̩o7�� � V�̩��S��75��M]4٥ջ���²m�!��AO��.�e�LeHkz�<�X|²g�ϓ�����@�'YR�w�o)�
ì+'�P���
{����`�Y:ʐ�kS�'����~��hm�jۆ�9�rVLeHr�
y�X,�����ԇ�Z ���0��2����z�� ��+���T��ֈ)�����:�VN��2�
~@�3��<�Ɍ�wZ ��+�V?o�g���ru�=]s�u������v��W){V7c��.��71�oM�v^���U�N�2�
q�X,�eHe�c�S��VO2�>����_�^����f�AO�+7����<ʐ��`�Y=��o��f�AN V²|ʐ�=�wKuwk�6����� � V�̩��S���� �Bd��!��S�`�9��Ad�T�;�S��XVO�{�NN�2�
|�X,O�R�̷\ � V8²y�!���&}R��ۓj�[u��u��d�*C٭S�
��go!�O2�9i<�X,Oq�w\�HfkD��J�VO2�9����
y�X,�eHw�h��;�|�1�d�*C- ��
��\�ַ�.�n�R�[ַ�Ad�T�;�S�	X|²~�3���C- ����d�*C=�>w�S+���eH}i3���p�X,�eHfkP13 ��WL�h�0RB�a�ȟk����2J"a�3��Aˊ�ƈH������.� J�s��k��\����>��O̩�AO���d�ƞ]+�8oWI��N�����h���+aY<ʐ�sj����X,O2�>��3�p���l���� V����LeHo��<�X|²{߯r�u!��S�
�`�|����ú3t�m�f�[5.���Y�V��͹ۙx�=n"vX4����9�U�1�٣l��5x�l�er�9~$����Y<ʐ��
{�Ϸ�:�`�q�!��S�a�k�rd�*C��S���d������ fkD��Xc
��� �}ɾS+��Ӕ����9>���[��Kf�Z���:�VN��2�
~@�=��� �y��NwZ ��+��������C- �P+���*C~���xAL@�8²y�!���?{�u��@��=��>@�7�6;j���b�~�|{���������d���:��kD�a�+'̩�}���
�`�I�T�~ֈ)�g߷�:�VO�Ri:�X{5�i�,�eHs��<�S���9�����IA`�m��O'Ri6�X)�|ʐ�����p���Xu�d�*C�H)���`�Y4ʐ�ֈ)��w���q�̩�AO V �Y7�����C3Z �P+aY<ʐϴ?&�j�ꎗ\����$� r9ӕ!ߵ�
{���a�+&�Ri:�
��ϸr'�R�AO VaY?{��ru!��S�
�`�q� ��w�
ba��̩/��D�1"1
cP�,��2bϮ����������D4()��r����@#FFy�C�nӄ"0BB ����V;3$(`jf�Q.���m<!a��u�t+�Z�]���`�
GU���l�X\�
g"6�E� ݺ�q�V:��6=�Q֎�*�ǟaw��qv�&�&]bk�*۫�ز�Ѷf�Hk#�M���-�8kQnƮH7Y<�nY��NyK��+�%KS&�#�͠�l��d�1�Q�u����?�sx�<i*T�V��Z��;���Nxh�<m���ic.�U��iq��>6W�"$�n�p�6��k�2Ԩ��
�1�.�cWk`̜�:���
SQ�`hōXV���p�,M2�?��h��@�?��޻�<ʐ��`�Y7�y�'R��>@�1�d�*C���x)���d�*Cﵢ
{��������T�ZAN�V�m���Y�k2�Ω� s�9I��N@<�Xu�d�����Ԇ[)�
�`�u�!���{�)�
ì+'�RZAO{?}�����f�AO�+�s��6��T��������g����.R�*��=fkD�����*A����)�
�`�y�!�u�
{�\�xXc
��+e���Xz�>� �y�!��D�a����a�ԆZAM�V��T����Z���t�����M��[�
y��
���>��������X,�eHfkD��Xge�8��T�� ��+�ɚ���u!��S��0���T������@�'�Rwi��އ��43�e�ku��I����d��!��S�`���y�R޴AO VB����^N�2�
u�X,�eHo�g-� � VaY<ʐ��
gs�xX,M2�35�
|�Pm�gn͚��.�n�աs�Ϧ�ɶ�7:�-<n�E�] �X�f���M�t�m�f��}eHr�
y�X,����:��kD����̩f��u�
y�X,�eHw�h����<���+'YRi>@�2�;�Ad�T���S���+'���4�Wmn�k[]�kw�����@�'YR�w��1�V*����#_��!)_������$f$�Ji�`�$`��u$���K�wwwF�5κ�`��` b�m�H��²q�!�H)�����:�`�u�!�ֈ)�
�7ˎ��O2�7i<�X,O��a�Ԇf�Aa? V²y�!ݽ����WF裻����
�`�y�!�u�
s3?^�²q�!��S�a˙����T�9�I<�X|²{?f�y:��H)�
�`�u�!������@�:²y�!�����ɧZӹh����'YR��@S�a���|�d�*C��S���d�����ԇ�Z ��
�VO�R}ϴo��`�Y<ʁ9��AOw�?^�²u�!��S�a��;�n�+˗b�f���NRr{�Ӑ'I%a����Ǔ����@�'̬�ߵ����a��̩� �=�~xX,M��=��? V��Ì�eHr�
y�^@�'/ݞ�׍e\�y��]l����{Sh��X�S�i)��Wg�{Z�ΫY�(����u��%WU_9�9?~�r�$���B�~eHg�w�xAL@�'�����ʾ$�a����/t^Bfܻb�Tz�O�64� Ț�F�R�8x�%�/y>��u��<O�½p�g�U���$&^B�} �T�D�ҪSD�R�(�`Ǘ)�p������/	���b��n�[�y-$BfW��I�I��M(�(�\!H���v�M;��_��0�	�U����O������_�~��VL��qAQ50L�BbJ�ż������B��.�y	��26��e�y#EgvJd�&t��#��_�q���9H��<mښL�L;�x���߬}ꛨ�ŧ��0��`�9%���DE��P���Ӻ6�h�j�#�k\�/v�ˉ�fCCB�Is\�+]`�]GK,U�.lgNt�ʛ��V��+iיL/v��%���}�(f
�H�虉&"*�"j*(�P�/�4�V���P�����g��ei�.�}�>�g{�_G~���'
�/��
f!N�~�2���>����^N>u�U���XI��Y�q��	)�D$6E7Z���䡝_Oԡ3̫��sl��-ܦ�}u����J*W�q ���R;t��F�fQ!��I��K˒D;��(a&$�b���t��h̔�H��s/?'�K���ն�vlR*��L�Y��v�~��_w�䣺�
e�����z�`�,u�)��.$������X*�.v,�EY�i�W��ˆ��M�����Z���T�x۞dz�n{ewM:�)U
�j3�8XQ�&MB�9�ب��;qU����Xυ����c�X:d��8�.$�F�G�
r��{�4��_T��3.���l���Պ��F)����{m�Ӎ�T_
�X�6XJҍ0[cy7�;�$��i�WE2D�w[��p�g�ͺ���D� �&���i���$��k���Ƹ��2��_�୊�r��_F�w�ӧ�OIy߽�9�Ġ�y��+���X�\����|[�Vq�dD��?q�C�γ)�����nlP��5�p��6eC�x���Y�O�H,��h/!�|R��h�
l��,#
^Qc��&��ܐ3�d�=\��'F��a;�2�gN���CA�V�ȷ��O�}��xiMX�)�c�4F��_+�Nhm��Y�� �<��ɏ]���z�oy�G�z� ��a��`Az<q�y��1������߼p�q ��w�g����٭''�9]˫L���ދޓr�+�5�]�D�K�"@�_��7���fE�3�I޲|J�ct6r6�q3�	����Ǽ��@�#��f/��Lc4�#E�O��c����砏�L��8�p�X0��q�Z>򙱧�BA0���Lx�:�bmf1��!��H���X��rH����r%��<tix���ې�a��;p�/Q����J~�]]}TRl[� qB�#���"ɖ#|��+�R׹!E�م�q32H�b�g1�;4hI���Ĭ��`�Q�7�"�yL�:�q�c�ј6aa�נ���"ky���]��w��Ղ�S��0L��,Sǃ^_x�=<���/C���{���"*a��tvɓ	��ŉ��;���&oE�f}ٚ5�p>��=<Y$��,�c��Vm�'���]#��<���{�ڲ�'+K�/0�r|G��}8����s�~r��ڹ<�\d}�fG~�3~�n�#�Z��3�p>ѹ!DC���3�{�%�Kg}．��KOw�|��q8g�X�_?�yF&\���)����C˧��}�UUUUUUUUUUU�֕
*4J�2�\:��m�W6�;a�X�ku����-�����+�j�3��6k�u΃���n.ool�y:�us��nB��q�zW ����ر3��ft�1pѴc˝5v�i�N�(�����䶀TJQj�hU�WX�E�AdL�E����g�l^��ɜ�Gp��<��7�V��L똷o'�ں��w�K����/�cH���J����4j3�7`�0�mv��B�9���r:��V�����v��K8 ���F:`��skYe�V��q�gF֑�ϡ�����A�g�^���׫kvݨ�n��}Z(���͈�c9�Ӎ��u��X���'FG�X՞�4�`5Fmۉ�A�'kl�^�.�8��f����l���O�J��E@�\��6ݹ�|�L>B+eHM
�����B��٫^n=��6%Җ~������w;��ծ��Gc�����:���wbvy��x���u���y���]��ڞC�-n��`��b�7�C����l���l�1���㎤����фIf˶
���͘d4˒�9��wge�ۑ*+d��k�Zvt	xob�^�;8{+��vv��v䷔�my����ݩu�nݞ�'r�����qםns厔s�ueֺR��pr4�/�h�@i�&��D��6+!�Wj����)���D��[�wfpp�86z�BZyƶ1;�0 +s۴��5��9\Q,ز�f��k�ܴl�����Ϋh�U���i�xyD�:G1R��"��c	2��Y��#IKn�q�6ㆣN�%��g��O\��@[w�Z}�7d�=z��#%�gê�y97�+ڃZMt�P!�-��׋n]����+��l=x�m3'l q��;�������&Iٞ�+E��Ut��u=ˬݖ`ݤ{An��X�li��Mk�WGF�V?\��隸.�vf��g�v��
�k��Rؕ5p��N�'aܫ	��j��Y�;�`T8C��r<��7���:Z�wf��BMsƫgz��U�v��C-6�C@�����������s^��<���C�Bab���g[\LG�qr:[+���Lr8p�%&I�r�7��p	��A		���1 �Q�d!��$A�cd���� �o=URXSk��a:�Lʶ6â���8����
��%fi��������Ɲo��spS R=���V�j��\kq�Go�v[NŌ�s�ӶZ0I�H-Ȓ��ry-��e�%R���3�(JK�� @ք��n��ě��%͞�&y�F7��#'v2C���EAmrmo�"��y�ٚ�wv��nk��V���n�ku��7�mV����#d��%'t>zq͗[re_�wwzM���lE��"�$�]$B�7y�8.��h3�wE�z�����s�w��ʮ�aDURe\.0��VŇ����L�Y�	�<����}�"�%�&x���Ѩ�h�D��,ꆚxƮ�//%�g�
�+�N©�^d�-0�;9H������6��qHK,F!M�JiqC0_o}�~��X7suY�����sα_t,8��b�)i�.�N�_ʪ�Ff<L̹<�������������.�2���-��a�9əZY�y{��Ц����wB�oQ2Z�A4�UU5R2E��m5z�Xώ^��]�U&y�����ك�RZU������S���v��\f��2������c�Ѯi�qrz\�K��3�x�2Vsq��ٵ)�j3�G���!2�0Nu�_��
�:�I$��=ϕd_t,8�ͩ�kQ�[�&Z�(�C��sP�}�2��!4��� B�$H9]�ffh���`�fP��B#bL�"c�t�ˎ��$EX�ip	#�i�;���S�_ӽ�lVz��.%3�^�Y�W˯�"|�eAH�N<�����d�#���M^�Y�{�J8f_D�y�p����:O㳾�(	�.`XJ�͟Y���y(���|*=C�u5J4�n���N>��A��滻��k�Z��XIO�'Z��t�Z����;���|�����|Y��}S����\���*9��I9��O�n�VF1�,s
����ɹ�
��e�:�U��ʪ�΍��98�b�i���R�,C-�?	��={�O9��|1�ҦX�󍶯����t�8����N���c����Z#'�$b���=�$��̔�3_d+�Y�>�ֈZY�	�6_��^�Sо!�$ϐe?�)dpJY��Zp�a��{���W�Q4d�$c��4Lp��]!ɖi	d�ER&�Q�W3ܮ\�)]s!�����q�B|v�7Ŝ,t�igǧw�:
43�Y�_:OI��D�����Be��=˞/�k���WJ��?(d�!O��7�N���6�ۭ�cM�Kp����<^!��S�"� ��`��-"aic}�*ج���6��L'��'&��Y��ѳD̴�����xm�����XëIO	��v�|��ʗ#����ے!JiL�UU�;�`��'K���Uk�c0N�Ȯ�Iyy��'n;�<?��N���R��-�]><l����V���^E�º�L��/������S���\��䐁�y����i�U���_�C�黹!��u\֭�rK�K�`���̻��>�奱ağv�4��-IvBk��Y�>��Ȓ�����~��,�YZP����k\+~>H �L�JiA����qwv:��QHJK�S`JhȔd����Cb������E2?kT"���c��f��?���R`��%���d�V-yt�wL�伔k���Y�;2��L�g����Y������|�kj$��E�RԹ��sp�A�4i���[�b�usK��WC��vKv��a!JTIQ5,L��u��/�iR�"���~����!&^8���ˉ��z��߾T�Db�F�uO:D���F�䗗��|-}�7�;�a���4�i��S��2���^�.�۽[�[6��Ug��w3�[0b�۩bd\r^��ό�|��G���B�ZQ�
>k!�u�ɭiV�n��M>����f�P�<��շ|UԴ-=�{����H������0u�	N0��!i��2��}:�-�Q��/m���\X�Ow�~��V-�eib������a�	�m������$���L&F`�)�b0�ww/+������S���Tn�e���,lɝ)2�դ����[FI.�����}���]���{�:��9���[�p���DZ�F�m�g���[F�[%q��خ�eH�a�>-��O�yl��:�:��.���M���Ri6vN�q�ӛ]]I��c��]q8�?�~�3�6����<q�ki��I�T�e&�`�jš�b
��
��]+G9X��lA�����:��05Ț<ݱ����{����wM������m=�W��j�nv��L㉣3�L���L�J���͆jCͥ����a�>?ۭ�I��������1ar���y8���6_����Oކ2�A
B�)���A)�i��]�Ů����;�a�UҦX��yV�+�K��L�/$�ϲ�����,�3n7��~'����L��V�|��Q���T�C0Os�g�mC���Q�Ӆ��s
r7K"�{�IG�M�_�}
�0W7ޥ������>�f��$�;�~*�2�;���ET*�n�&T�N$�w�g�|z~���t�B�H��IS��i�M^�X3��9'7��ߣ������YZ�F�峱���r\���í��0Mn�%�Uv1��	X��\#�QRR6)���~���)�Hî�����}�<�}䗺Ǿ6���L���+��R�[��j�ܞs�{�������LD�}:45wrG����L0IHc
50у!JX��H��T�=uX�*1L$&�i��>湙N���yP�������][;�{�/��r.�R�f�Sg��������>t�O�_��(��y8�Z�rU��а�*\ƒ?E)��p$�h��ΨC}�^�ew��̬�_>�-�1|-qYJ�Zr^�G|�|_
�Y󸞩�"I�����E9$p��;��ϰ�C߾|��\���o_X��_�fF\R��fB�{˿����w�EnF+'�$�1��[(�\�z�jw);v�uĺ��iVe#FPBPCs
�L����,�|S��ZEB�ݷ6�g�����{�XυM�a~����Kރ[\)[3��_�O�}���K�q���T��fB�y�[,`�:͟q�> f�N���TA��$n4 ��F~#�}:Đ�"{���bL*I021�e,4KݸBI_��4L��EI�fX���M��ף@�����^O�1OW�ZH����sm����<:�OssYY�p"�>9����ϡ;OŜ,�t�uL6w�V�l���\1ތv��oߊ�-�3kwj��	��������ib�r^�Z���aƕu<��i�
kuŲ�,;���o���H`W��lܫe�*��>fS�;5�V�{jՑ�6w3��98�"�;�� -��H$_~)�N��ߞ��C�nT�-,�����I!`����e�*~~��28���a' �-CM>4�N���(�/�O��N�8w	�P���kV����G�v�>�Q3�
*D54Be��Eo8W�5����u,����y��}� �ȕ����_Y6TD��T��U��r^G�dY��.0�_[�v���4Z� )��s&�c"gv�I��h4H�����n�e�Q��ڈV
��Q�)���Ͼ94�Y�]�ߴ�iF�K
���|s�\���r���1�D�y����Ϋd�VFۯiSK9/)�a��GEMx��6f�6��\���i�v�MZY��K��h60M0�IF�*�e�Z��ݗ���=>��j$���`�nϋ���X�]�r��?u�5���x�:nn Ӊ���ĉ5���p���[�Y��\��3	�t����G�n�UBӗ���C��)� !#�>��C�#4�8��n
�����|gEGĮ≮N�3��c'�~'}�����Y�yg߹$����£�H��ZQ�
���Mw����y�a��?S����+r�sB*j��V3�)3�U�/$7�u_p�e�O�sL>�o�Ň�JxB�w&&4"bjH�)wm�;D��0 �tLĘ��7#O��n]ݯB^���e�X��������驭�e�HSFf�F��l�y��vzY��b'f�jy���z@gm]��`&up�!��C�K�O`��ez�i�Qo��T��6�(�Ra1��{��U�ֱ�#5�X�×E.��))��;z{//4�^"x�x�1:璡5�y��w�ƛ���4v9Ӕ�18�{;�t�r�] V�w%�#3�����]�&$c�]A�jn8�d��ۮ�.Kt�e$?��s��N/�ܶ6ƧN�Yp,ƕm�J�t���F��7obr����K�X�c%���Se[�l�xt������A�]�V�-=��R��O�|q�S�BE?S����IԒ)�ß8�E������g{�.S>�ʾ�vڪ�~x�z���|��$�̧[����ɷW@�!	�"�����j�P�N5t�ǻ��>�W��Ŝ/�S�i3L>���ʕP�Ңi	��-���x�s�SI�3{�Q�����i�^Bn�x��_|P�X*�Q3Q34Q)�Ҳ�?�[0b���ݕ�MBf��VŇ����L�L{˸���>'��e��c�7hܖ��C����]�f��ö�n�o�8K�ٍ��l�.,ڋ���P��MuR4�i���޸T3�/[�G������fǮ']��o��YNU��QT�.�if�ܲ�i�Ǔwk�� \�wn9nÛ��0CLM���*K��� Ɠrڂ� �$����3XZc��U\���p� ��ӽ�P���G�")����D��t,8�da+OiwX��m�w��}I�0�d=�b��L�}��C�9֬ŝ<>�9%�#g��~��/�qq,�i��u��� *��<��~�qq~�"RJ$�MT[,b��7r����rJ3^t+�Y�;����(���8�Y���+�";:�,�A�FZؼ�R����m:͋5���!s:��j�,`5RS55֚��kL�T~,\y���
���g�<��Z{K�[���y.���.x\D�f��'���%iǔ�?i��H_���|&�/b�gt+�wS�O6�����N_�Ǔ�~��R�A�����Ξ�G�}��i����,��7b!6��H���u�����m4��-!�M�{0Nrg��޳�a��{4b�XG�V�)����'�͟ã.7/������#ob$E�^#RMN�C)�kO�/�X�p70��:����|�$#�j�p�[�#o;T�c�IqԚ��ɯ���H<:0�w%��lNL�E�D�D[�xF&a׏9��}ً�/�H��G��܏
��W��-�U��H�̎�A��n��1^{��.�*͙�1���;3|w�ô��,q/�iH{���in��u<$�����k47�J7X$�(�Gt�X����ґDՅ�}|��;E��S(��X{��A�����KI'{�ݷ���Ò^LiEB�D}�,�󫱱Vpg���v½$Sv1�}���I����(žs��a�IK�s۱�_Ez74kZ�'<�L�<��ܟ4�͍d!{ۨ{PQ"#�q0�y�-5D�Y!��3{�:�nk�!o�����\Y��?�8�1n�#`����$���ɤ���B�|r��ܟ�v��/���W�?��]�3�s�g�OAG���?!	�*y�z�V�؊��϶�(׍f��^�kc=n�d�jb�)��33��|߷�[Vso�K3����Vn�n�0���\K���Ys���C2�0ͫbP��L�l="3'�+�s���4�ymZPoDŏhmgl<	�X�<��lM�;�x{>�O�/<���ޙ��~m$�7˳y��u89��2�3����7�^Ӗ����dU���c}�Q4�h�$��YB`�cw]�9\�.�$/ڧ�����^9�3��~��6)��H]���IB��UD�T�ҿA�;�
��)�&y�C���X�"��i�;�Y���}W�,%m�GY��pe�eӥl������,=Gyy��TJ��`�럋���Yj́��8���._�C
�D��MC��X�[Yk�v�&��@u6��e�,�L�s:�̭u�6��l6ڻ��g��g����ʑi�2�=y�[,b����w��p����p���6�̑PU��"��UJ4�G���\��B���Iŉ���d+��[��%i��B�|���s�fUv�6w��O��{^��[>0��qlU�^�|u�uA+�����A�l��_3`�r�Z�J��I��/G�ge[�Vq��-=�d/��V��dc@�V6H�db�R�`Pb���Lb�A�]ݸ����c"�����1�)�u����6G���P�!���n�<t��"��+��|)(Z{hn��±��'���=��s:[5b]`�8��E{R�v��ۇfۑՊ�]tFb�,f�`�\ڈ���a8�,4��
~�u
?f��K4�#f�-"�ig��&�{�|{���%2�i߱�JQ) 2O�P4���x��S9/T&{o�����Ɩ:ȕ��ˁ=o�S��q�Z�g�Q�"�B��̪��7��+b��7n��iG$�|(������VoE��,Zz[D;@�)7!q� rB3�o�>^?�,�b���	����0b���+H�Zw��2��|$��C��8scCr͍����57�ߤ�
��G_NR�(L�u���c>9�KOiW
�B @ c5����2K�d�1PE#d�%r{���
I4V�ߟ���ob��0&^l�&���U��R��}.��m��n��f�6�e�_$�^������D�&7<&���V:N�]�ē�C��蓅�WŎ�O!�f:8� ��n��q��� ���sƷiqq��`C�@���J��F83)��g�+ѭXn��і��qY��^�u���sZ�؜J�T�rו�3��C	�u;��&�u� �[�����y���,KrD�p4Ě���{<2��:3�n%U�0�:�2��z/#{'c2�YnVX�.��'������WK/��V�g���D��2�|.����Y��K�(�3MX�����Z��n;�G��9Y)�fd-�ql���n���u)�o[�	"jj����~��PP㇎��՟Y�'Ҿ8����D�K�sz�P�TΖ�d8ZiHQ2H���~�/j-���G(�	�0������Y�K!u���������������Qm��\+���X�\�u�ž��_,��i�/!n�?�ك�/"�NAUT�F 7X��Sj�n�����ِշm�ncN�_^��i��b�"iv��؄p-s�!J�S���R!�K�ؚ��H�R��䐰}���Bg�m��Q��k�#��ݱ:zt��}yhC��$"5���y{I�B�CI2�@3d�#L���lߏ�!|���]C"�i�^������������Yh��ѹ���t�����~�\+ �d�G$3�wW�o�a��^���� ��Z
B���$[H�U6�{���O�S	�9����>�PBҏ��к��W�;�Y.����U&ˉ"	n3����kΨCO�d{�ed*���C�k��L-0�������ΈL�ˍn����ܠ�h�vk����LX���6�f�5��յpۢ���r6�q�D?Cn~�!N:B�Z3�������t`��}Y*��|q��Ù�����D�q���3P��|���F-E}	�p�e��-��a:�T�/�������_��45��&]����tE9�$Z{a��n�^���.[�ı0$�(��B�a�������H��m�/�2��3���H�*UI 	�P!��_S1��o�:��T>D&Y�
�m���qƊ{�+�=.vc�)�^��
Q2ME�
�iR��B��e�{��f����s�KK�ZY�_:�,=g.���J&;u[n� 6�x�/�2�{Tz�H7u]�\-�ŻN�ia���9��Ƙ��.�իɕŌ�l�8�X�,�l�X��Ʒ�Ҭ�=9��2�u�� "�Mz
��-�1|Q�����3�<�|+=bݶ���i��q�߻��i��D�*���~�XER�,\{O`��_�E5�-=���'�'�����;���8��KY.�N�r�)G�+�&�3R��_���su���4؎t�u�h5� �F��XѠԬUE�����s|��Ɵ��A��`��q��jݮ-�1g/C;��qw	�<}8[��|���x��r��?�%��a�68�tH��� 1o=b�kM�q�����vmZ1��XU��ui^l���)��
%�$Zzum9�p�f�YU�����:���������Z,��E�I�0���l�#��7ީ\X�k�!_�n]��p��I
"I�pD!Iŗ��<r�FG��-��eд��8L���!��V�G�m[����@�a��N98{�^#��y�}�z.�t�i�᜶3�ȠL�3!O���(�"Q3P �I��d�_�pL����w_9����ʙZY�lד~��_����(�̕�[�$�$��Dh�Q�����u�J����U�8RgT��v�fd��I��E�N>�eM;ng��v��T�T��W�`S��l�peE]�ugml��Ǝx�<�	R�[+6n�J\R̭��Փ�ғ�������@8�KZ�����u�ԷY�W�\iʾ�8KL�u������\��a��6ẟ�v_�/܉�V��=n<a�d��u\����͹룞w8����
<�Ǆ�>]*� �3R�K�r4q?�*�g���A���ތ嗴k,��q��z�,����q�w�GjElJ�1�#���ffi�g_�����um���@�"V�Ү�x��{����X�g��Ξ��[M��j�e�(���a?Ch��,g¾w��#�_
[��(Zzu������s�ԪT)��2�lS�9�p���)������q��M���8����0U�sZMS6�$��g�m_����ǦR��}]�^�_ѓyT���y*��b�O��;ؗc{�E�L�|-�k{����Y�]�SI�3����i�;,�?~���ȓHђ7�᮱�\�j�q�/u�hCS,�e�l�Z� �6����+�����r{���E}�
�����C�-�1|S�b�p���3�y��u��N>͎�ZW[ߟW������}>~w�D��%� �14���h،���`:���t���>��͔�=�n��±��ʥ�	���o����E�hS%MM�qN<˘Za�S~�,�G�+c��i�?g�>g�_BZtF�s�MQ3U��yG�{�V�iW�����C���)���[�9�q��q>q��%70 �)~���~hS�����W�;�Y�6N�-=:���C4������T,���5B���k�ɗo:��x������dM<8�����n�`����$��O������S���;`L��͋q|��}}SP���.���kp����I-�3�6���yڃ=���W��,u��i�2�m�K-�ۉ���kIh��ͪ*�[�c�S͗�}6�g����S(��@�����Թ�TDh��c27KtNk���A��#-ѧ>g�5��0�?t�F�)Dp&�Q'Z�7���}�S�9��o9[,b���=��-;��||_
�`�.���&����TU-,��X��f�Y�B����t^�T3�Lw�)���?}�G�IBR
�a):�gV�nn���[Z;Mv�s�w?�>yk,��V큤�����J\������=?����P��>ߜ[��뜥3�`υ��߹�<?~��s��-����3,Z{�/n8ӏ�ȮP��fB�}���Gp��w)��������E"b��*���h��Re`�k_���_�7Qŉ���.�����
h
����$�54�������ݴ��8_-״����ȶ*<x@�$�~�yW�2be	�R*�ej1V�^35������U��PL�k��&b���cT��B�rC��*��a���T�������6��8�|�BSQ"��0c<��m�6s�iMW5�&�L�� �K�fd*�5�c.��[r�)�[j���X�/{��g��[���`����T~���_�b��)����D�_4[���gT0��]kJ~㘇N�NS�����*�if�=�b��R;��R���(&�	��:G�j�s�6���%q�r��W��.c���iY�o���.u�\m3�Θ�?����:-Z`�=�lTz�6ڪZY�
>�q~��4���w�iB�$�1��p�~�[p������≮N�w�l���Wv/ㇾ��0����>@w�xP���j�)x;��ӛ���ԧ�!~.�>'�7�ֺ�~�H�}��y�!Q%I�f��G��xRz�N��m p=z���ֳS��	��򜐾��`�1!4_�B	g'�=��z����x撶�d#���.����فfj���Z~\>�Ha偉�Dx4��ĉ��	W#��Y�c�&�����'�佲=�ug�}���Zw7L�LK&�Ͻ&<l�V\�l����'�ذ�Gpa.�D�$:ڋ�١9�{��q�T��?b�]��݉��LX^����h0Cm�d0�8Fyl͋����׳�s��>�0��h�ޓ'�!iYf�!��Q9�-I���C&l�����]�M1�'��`N�F~������;'c�B1�b%�/���� #����o�J���?��џ>�35��h�<��������=}��V�A�<T$�+�X�!,L넉FA�6��aV/���ώ������ۭ'�Z�X�3qy�\��T7}:�(�猞����k���N��A9=�>��w��Wg�k�C}��FN�x5�c25G���Y�c q)+f[�nAw��ûv�=��`:QFH[�/&�x4ǔ�n��S"L��FC�ƠH�4��{��O}�~7��RW�_�A~��8o7&&'�4�?*�����������ֳr����Ūۥ�Y`,�k�:��2F�ׯ=�x�r��&n7=A�%L�=e6�e�.���2�i�1���t�KŲ��Z�8+�5��� D��K�gs��]��e��7"�m6g<�s��;%�q�#��si�y{xm��S�U�.�@w6z��*��m�rM�9��sB�(�.C/��N��r�bg���Œ{>z��ǘ4rRy9�E4��.vm͆;cÁ���F���pm�3E�1����:������]���l���]�[���&q�Dǳ�� �UY��܎�ݸG��v��\�"���Α��DX�.��� ]�on�s�n�kӮ����2;J*���Z͸�j�8h���ـr�М�㫅��.���a�ٶ"��%���ظ�8��1�%C�{e,��j�dw$��6{ � ��8�Q����[RƷ9dc�8sM�䞛o^Q��=F�Y����6K�($w4Jk�DbL'Z3��7
�"�E����^rl^�7(����s5k��a��L��ڑŸun�/\j�=;.JDz(9�xn��!-����+1RZk6��ChV�`{��.��"�	�%�u�J�1,\p�H�],�֣�z:���X	�*��a��˦b��f*ض�j�Ma�F�=g�Z��g�c�{L6������2����m���;��`����^ٛky���#43Nk+��O7nB7H�cnɶ�g�ܭ�lZ�K��d3�s�@ع�.zW�'Y�t��Ӷ�D�����l�K�M5�w�5�#Ȗ�bƛlv�r�oF, "���3x���'8�R�+�1���ێ��I�\�]�C���p٧�:�/���-8�	th�zR��/��n7�5�<v�ո���9Ψ˖筩���� �!���2\Us�\��#r����ĩ���Ѣ�F���3�Gx�H�X�`]g�Ds��k��%�-ly�RYci��e2�
��e�K�vl-�vjX���5�.�v�]Z&�9ݮ����*A���(��b2��$�y�׀0M<v�&4Y�����"n6�rMu�niF�3�N!�+v rc�8�QEM��s��ݔhƤ���DX��HrR�'��=Uf�`�vX��Ms�C�+J��A7-�Z-1��.�k���h�tR��I��M'(�Ȧ�&�m�����<\@�Σ��#��+3�jT2JQm�)E��[M.e\�F6g�n{wT��i��,�O[]s9/��:h�=����B1�]1Sk
[�
��fIu�M�5�؛�h��+�����keJ�f�G�	�+���F�vrٜh#�ؚ�sds�V	獛+G��#�^�����n�2��]��ĝ�|��;�[/f����`�5��o�;��x{	��*!2�0U�����t9��Iŉ�n���|q���Ԋ*��"TU�URg�������0�|>�_Be�&Yod+b��}M�D-;!�
-hC��M')��?�!�9�3����w��}E���fBks��f<�YD ��b(��f!߂�m��a��}$�Y�	뿡_���?yo���Ӈ����h��M���W�����-=�dw���b�Åe��c��q��^�)��jEFH1Al5q���,�<l�u։D�pE�!���](�6��͌�K�t%y�]����L��*�cp�u�t�i�ٗϥ|q�L_z≮SG��DR�m��t��<�|���	 �ry����@�	�4DbA�A�*�S4���|*=�u�(�[N~�дP�J�i+3��+��'N}_�>w�xt�͵I��8�!k�پ0�X�N���n��S(���F�_B��)��Ǳw.,f�{���e��I����[�Tq��ș$��IH�D�Jg�˅��sl���(��+̻��7��-�Y�n�P��Ly���j"�b"��'�;��f3��l�V�sZ���de�E��]�[�W=0��s��ki�m��Q�:���ŧ��e�
�iN+&y�>�S[ܯ�8X;��@*�L�I%TUT��P��[ܥl�a�+zzL��-��*�cp��s:vBg�B�uT� �+�(QM
��a�+&�i�2�~��k�x��E�PTE��XQ�� I1�x.�R<�2�0���lT{	>��fBQ�BԊ1N������gt,9T;�҅��V�m¡�'�y�����[�)�.v�w�0Ń���K�Z_FWr��R{	�|�L�Lu�o�7
��Srt�R���*�� ��fJ�����l�������8��n�,D
��mt�u>�cw���-�T3��d�)����x��{��v\�U�f�]�q�AJ��QQUlXz��䪔�0g�֫���аc��L�i���W��W��,jN@n8��1-�)f���� d�w�|Gw8W£�2��Re`�����(�d���H3�=P��\.�#O=�~��`τ�.U-=�! 	 uJ)m�6_�I��V
"�1R �{�B����i;�z��g⩩ha�Ӆ4������,��!���j���:GZ��>��0�^I~|s�v�Ţ�l�J��m�^\FVܢ;a�r��˧��8��n�ahv��p�1���2�N"Ӑo��i�|ܐq�/!}w��`��ɸb�ѕ	�^��y����;޸3-�5GP�0����&��6���:�,�3������d�)����Ц�ܧ���"d��D�D��p�ח^���};�bΏ`�)�*W3�r���cp���t�L�D��q'����/�/�Y!���WS�Z{K�T��-�1|Q��ZMBӧ�^�HT)8R��pÔ�?i�����4�m�u~��_�ԚP��c>~u��MK� DU��l�1X�dG��U��k���{��Z�m+������G��ĳ�j;{�7)pl	�x�[�-Vȶ��j��XVj�]
ܣ�q��͓N����G��#�]�dwl6L��&#���Wt%����-s�)������+�.�<��؊���s�Mv�q�ee�6N�6#��[lܮ�j���ʭ���R�4����3n�f�kl�K���[kq�=�<�󷧴fܓo&� {hq5�@�`�;\-u����.�'�x�y�.�{$rg��=;k��7kl�*%W��s5f}��ιݬ���g��MJ���*�32��+N�5�ബC��Ӕ�~��^�㇎��OZ��;�,���1���w\t����޸V3M�Rg����[j����#��ha�G�V$�>Y���o�
ذ��V����7�*z�zp�����zI(2Be&S܄=�8����We�.��Z1��n��M��w^yH��/˓R�n ��*��4�=_�nw6V�-=?;FZ��x̎�)��jupƣ���n2\N�,rN�M
2�@��$F�Z��m���΋��ɑY�m������Z���D8�]}X�C?Cj�$��/v՟CjE6<����&}�pk'��9�N~�6b����s㠱b1F M��_����,ŵ�B�̬�[���,b��W��t�J$��1�
	&��+=��k�S(�[N~��t�:�'�8�3�sȶ�X�U��DMB�T��!��S��-���a͟q���}:�-�u���"3�7��h$����g�چ�Q8�8�{��m���;ɛ!3�^B��sl��
�g��Z�M1�����\ז]�c��Χ���.��1�rmn�a�ݫ�'<� m҆B
��3��=^R4�����b�i���������ib�����	*$L�,�x��/ྦྷ�
������F��iUL��V�ھ������S�����pD)�N������|k���,�HB	( �E]�����7H�#���-�/�4�{)��.��5'�"�RL@�&S?�������Lóo��Q�'�腥`���O9N���t{|�e5��]�酧�n�^�_Ӻ>�*�e�&�:��im܀S1:z����P��0?���yѹՇ�7X�N8��첓�7��KW�ۙP���31M��D6I��xs�}�	�i������|&��'&zm��g��i�x��-���-�Q��q1��9�Y�FR�#�,q��t��H��uz�b�<t��	XȬ��)h�ϰ�C72	�����r�>��N}T��]�e�F,����q��m8ԋ�[C�/���?�^�UD&Y�wU��qH xG��o��ݮ�!%#@$R��y�*p�?0���&0��8 r$�#:��N�Y�Pq��bξX����iWL��lTz�� ����no`�d1rM���u�lz��n�9�HQf�\:؁�5��;Xv1Y��ب��Hq����:��3jl��T�8�T�2�!�H�5���3�툶����IRL�M#M���Nbt�k�[��h���`���_�nǜ�p�qFLM��4�~7�ӝP�N���(S��[��H�'K)��Ӿ�u�iL9����|�<9�����:G�i�>�jmJbt�~~�uCM<s�R��$m"ےH�����4��d�Y�c;!q5	�C��V�G�m�MBe�`�BA�r�y%��b�wwl���>���6s�69r�4.�S:���k��mL�k#�Tk�b�m��j�s	�֘hݜ��g�gm:�܁�Η��lx�k�nrT��-�Aj@�6`��1�&�-l�lQ�9
�j@��5�G`�"��w:<���y��j<G��r{Y1��Ų<7%y�=�*�e�:l�8�N\�p�ki�9.-m��:����ƛL��,�A�[��EtՅt��l"��2���a�:����g@n�a�t��U�4���8��cVta2��[6sP�&�Q�j2B�(��4Tr�������.8G��-ŷ�
��3�e���l���TUM�W�荂_Ĺ>��t喛g{����C0Z���Y��i�G���0�`�!"ӓ-B�|'�sKOi�	��M���X>��&U�e��lV{�Z
f�%���IB�<t�ӫϙ�]������q��4�6@G��!=��!n6�7!)ɔ�i܃��q�lXz�طꕥ�`�K�7������߷c/�e�	tEqn]�W�m�f�\���I��{<3e��
F�q�-'���~�r�0��1J��9�Ko�S#�K`[C��vH�&�f��O:Lq>�t����GH�F��׺��/��Bw_t߬w7P��{6�m���c���+A
?�a!j8��u	��-�1|mӯiL/v������b�<t�2RR��� ��ϙ�ᩧTi"�Ʒ�m±�(�j�=�1v�yN�G�dpa�Jba(�EQ�]��ϳm¶,=���"e2�0U��ϙ�,���dq�֪�(�D]���[�=b�ظ��>5H&tĲ�#;jm˶�*�=[�]iJܫۭ��u4�A?q����e,�0�w 㘇>�y�#Oк��H5	�F7�S���ϰچ�dt�Y~�v�ꇍ<c�R��q	�dM� 2�i��9NG�=V��8��e#< &��Y�'�a��ό���Ase�l3X���A�2Y0�)E�l�W�D܋BE�q!��g>�x26	�FjO0��!�9��ݾ�5��{$�vvh��;^<;o�g�֬�x�pM���m���? �"5G�٧���/�xo`�Of����{�ݰ���Ӝ���?GV�`%�uH-7}���E����n>_�!��m�ׁٗ/����6�^��@��Ӵ�&�H�aF3�K��7ې�1i��E�<[�9`37&,���?4f��8��W&�{��є����d �K��v9��pC}���x�ǒ_v���#<�M��������h��;�#����/t�c�5& \P@�E�]9��Pɉ�U,F.9�䈁�y��֐>Hx�Ti�g�?c��f��x���qc3�Yy�A��n���,��F�-�̍��/f�#�OLE�N�&l v�<�P"�ǥ$��w�����_#�n>9��y����ѡ,�!�?,ƴo���{,��{�)�
o�f���p^���4��.�̛�]�T�\�`��}���W��G����Ŭ�
D��ʥ��{�Cs>x[�.�8�2�(�D�o0�"��Í��ĝ��I͚"��U��&#]	��`~�&��$��ݾo=�B;[�|��0���5���D�./.�~l�	�~�ut٤�RE(s�0H?�87"n�@A\�9����i*5���ї�u��hJ�͝U�4�}��7����P�A��T�UW芋�x�3�ݗ
ۅ�ϋ%�i�2�}{�-�1|Vӯ2*�[��wEɚ���վt��I���Y�:B�6���i�׍S��N�e�zt�I�w�.m��`,�b�jM�E���l�)9����3�<�멉GK�E"�, ����jB�@����C�o��i͟S��=e|r�о���x��c$��e	H��6��J'G�r���4Ӧ�SS��q3��c��w��m�e*�|-��r��Y��R��L�-��f�Xw�������{���TV��]z�X�,u�+Oi�
��e��/�5�/���_��i�?�^�vɠ��+��m�?�3y��ɶm��~i���BO�B7B�x���3�6����o���v�-Cƞ7R�Lq���l���6���K,!l���j������s��LV3[�)�]Zx;v�1M�#v�`1!$(M��t�<e���ty�b��KZ�ZQ�
�V��I��
���}�Aa�!�����(��`τ�2ii�.�=}��s0qƇ5�i)sE�NXe�R0��D�,�����N�+J�uxr�4��	cAM����mG~㺇\�2�iB�qq8cu������HL�L2��h��KhS�g�چ�V</���Gh��|3JqY2��+!M}��Pł/����`��=�����=�����3�Z�,v��-�ڥ��5�A�hř�ҨY���<rX��t�6z�-y�pcs�K�˗V�2�B�i�g-��%�f,cR�*�u��1��)n���n˽5p�`ǰ�ϑ�杪�'s�`�]���ɶ@y�=�65͋[ 8�<q$s^��ʁ)��Clp�zʻ�Ϭm�η��=s8�Q�[m��,�A�ӏ2F�:��n�����v|g�0�۩]tu��,�V���H����n��V.�q֗Nù���J� ^�.; h�9�\ݥ�I��Ξ��w���Ig��n��iF�-��U���a�������{��scy���}�<:zG�dR��e�������%iwK2�NR�M�47>�}1��N
�J4�F���c��H����Ӥ]�pS��'��SA��.@�lF��t�<zǧ�f!�{����?i~���0��-��CjW\NR0�a2Tn���Kr�4��R���2��-�1Y�˔ʸZ`����Q%[5Xff۩P�hX �k'�Jx�jϰS�q��w�.����+sX�N0��Z�e#�}U����Z/���چ�j�S����p�i��b��bPD`jnH����$�VS���s���y��C����t�#�).awB�f0��୊�xN�w�O�IS�K�n�*��W}�i�5N��.�NuCƟ,� ��3P�e�)�H�F��Z��2`d'��)�:r�Q��~���C�<t�x����P�D�CK#��Z�0������Z�4�7��5/��V��ɳ̻��e7�b��3������KI�����h�g<g^��.��Q��/O���5̹D!�f[��,�]���p�)��H�n���P�ly-<ml2�±��M�&{L�S��a��� -#"re0�4�� �0�{�lXzϜ[RJ��0_<x+����wn�t&k�s��*���|sV�m¡�P�"Sz!.��� �xB  �T�2�,ͅ]��(�|~�63ㇻ���"fH�N&L��#O�l�aB�x�����6����F�G�]�2�<iӀ�8�eF�I�`�%"q��jξYN�G��q9P����qlV{	�"S(�_��K�^�����F��k��"Z9q�V�hFh�������:F}���l��V����(�I����C$Zxm�^�V3f]Rg�̅�jك�18�U8�a���H��8���T2���>����4�S�����Q-���O}�c(,��a	EB��:�<UX��O�f!�o�S#L�T8Ƈ>������Ρ���s�\fVtO�A֯jϡ�4ِN8G���:���S�[���]5���DEr����T�<��.t�R�`�����8i?[�"x�=X�C?C�er0��;��ϰڇ�蘠���[�\��y�ֱuC��&��[,r��lw�ɮ/r=�A,-��6�������L���o_X�\/�|(��������ݣ)�H���J�8�C�����	ȓ�(��)~�����L<t�����P񬫍����q�T(P�H�hE�P`�c��s�f׃�ǌ#��x���Ӕ�~���	
a�Q_agb�T
�-��l�'^�����?k�
�|\ſBg�˅-���F���oȨR"�M8���C��_<-�Y�������`��?_�n�=��﯏/��I��u�K������%����U]��Yu,�n����ՑWi�NR�����E�G]�F�Ѡ�)�ͺ�|k��f��q�&{v��k��Xu��qo4>�{c1��Ԍ�6X#IJ)8�f��1iM3&W����PѮq:	��hL��qV��]]��!�M&�q�]�̾y�<��֫q���3õ��1ƻ/&�h�Έ݁�y'B;i�2؋��`̭Gk`xJ���v�y�]C���]�y�E�ͻ��/`qB���am��b�h<(�m(t�;#�˭Xx�S^�5��w3��3j�y������!i�/!W���e�_
�w+I�Za~�~�F����0[��nCx��vg�mC��2>8G�ٰgT4Ӥ)��8��bRJa2���82�4�T�St�VR�O��x�����mCǙ��>DD��)H�G��VZ�4�w$����o[0b��p�˘ZX�ۚKe�e�^VI�I��O���gǇ�
��e�F�|D�d�OO��녃><4<��9��Ͱ�b\d�jhq�	�.�Sj�,̈�����1��%ԋ)fv���6 E&�n|��� �mL4�#��&M����lX{��$���`��Զ���� Q�|��a���r�B,�W����w��������_aW�Z{K�Uz��0�<k8�HA�FY�2ۓ�"ai�nl2ب���T�&Y�u��a�6̐��8��(e��e0�2 ��gT<i�Q	~�5	�YNG��g�q��Nt���{�X�e�)��,�d)�a�N�g�ڇ�f:�G�w^uC:UY��?q�����f۲�Z��;JgMy�m*����P�O]�u���&[Xջ@IYF5r.��q0���(&j��1`˨be�-0���[���r����`�w�ߨn�숛֘�4q)[W?��oO;���z�)��b���H��.1K�8����c��P��0$�F����HZY�t��߬�� ���H�� ]�1Gu�;����|z~}qm����/;�Ʊ�7+\���Ǿٞ�V�����2��_�c-��`��[:x|zFG�"�Y��͸�|�p��wPiB�����+�C˅)�����)�H��e�ȤmG!#(�.-� ˞Zd��L+W1�8n��]TL�:gc9������[Fb�+�������e�Y�6�tL&Q�
��q~��_û�LO�Vv�ғl�l���o\,�/.�i�/!}��m�1|'7,�q��?u#)��Ph9S�9�8��
B�x�ݕg�ڇ�}p�a~/�C-B|q݈O�w�+���i"Jn,�F��\C�u=�b��|��I)�i�  ;a@��*E"�m�e�Of����s)�嵇���P6�Q�q�8G��:���.��&{L�R��-�1X��d&>Y��ߧ��]�A�e�m��K`��L�\]VSK��4d"����hs�Od�&BO�� �aڇ)~���R0��}:����±���e�O}[C/\/�i�YW�4��(Z.I!S��'�j�p�<g)P�D8��K�)~��VmgD������[X��\���s�i�׍S���(Ψa�Ɯܐq��j��e0�<eQ�J1$¤p�L�8�]M唈~��ؒ��\�V|ͨis�q��Po�@��G���-Bx�ְ�O�wP��C�[�ZM����ձa�/Ƕ���� ����4,�t�� �hv��!�5��`Lǘ�?f����Q-6O�0b!n�ձ��B3��	[4	� �B	1�n�k1IH������� �065h:�O���l��P{����׺�r����浣-��m�C]�}��������?kZ�fŜI~#w�,��;^�H�!�%�=��-o�$��/Rw2O^ףӥm����(�1��!�Y�����!�p;��g�g(`9'�[1?���b�}0�.1�B�&�
�m7<:`�(�|�����[����m&<8��3�!a����=��3Z��F#��#�^�|�Db��Ŝ�������
�����F�C*,8�����E�����Zq�	d���Sޛ<Qk��dz&�,�ug7��QѼ���V�D��%n�[iO��'�����D�F(XP����<�.I<�-z����OL�%��x���{���z3be`�� !֋$���8t|W��1o_x���|Pa}�$HlC�6!�~�E���L�^��7��O�6m�����*�􇯳���Ƿ��2�?6� ��1ב�����Fǖ�e~��e$֠�2Wa���z��{�3C�odHFs�Z�ڳ=�!����?�o3�pL�q"�8�C�6�J&A,j�e1U��m9<<�\�A��_{���d--,$���IO�{����7���¤�>sy�ʪ������������ъ8L9�vvk8�۞�v���L�8n{P�ݭ;���6� J��lǕ�T������A\�t�Sh�a�j�W���������6�b��'=��� F����z�1����t��X�y�l���>:��7���/YRֶ]�e��Q�Νjݸ��ehrnc�u�nníչ��]=�t�E;�nnm�$�n��p!]v���u�ؗ��V-�;������X�و�Y��:�#q�9֝�����OHg,��q�J�*��SX�6�J��d�k��$o\���MZ�v��d�ƪ؈�vlҼņ0�]%W
�4������L#�N��u�<x�<@#�6[���[�;�����m���iFуyܯl�u������nx��(�y�U�uc�yz��:�1Yq�(K-���h�S��t8t'���7meě�����#	S[��/�v��z����)���B��Z���N�E
v������k���W��l��Xq��ZR������,nc��v�+�G7Y�`-��m��T#���&ku��bM<G2�;�ۓ����Ss�Oi �nӛ�G��v�J�dl*g��I[=�.��{�&g5��ݸf:Bۖ��7%���t�j�c��,a�ɦ�3u6Yݫv�:H��Y��݌���
���vASc�5�z�nSٺm��ct���6�n���R���$�í�W�}����l��b23�.7[�-fn��˷��9d9n�f�x���j�pu^SZ��l�\B�6-e�Txj0�a��� Dk��^WY���r�(�h:'\�{��-���]Z��=N��rb�/��'4FyՖg.�ŧt�.{pP���}q�-�A8�N������'=�.�3.��i�Fk[XD��icap�P��ǘ�H�<�X��3�vI���	`Fi�w-#4�E�.���!!1���)وݞz̲.�[�IܛЯi�<ڨ�f�6ٳxKS3,v!������C�筦��v�G��η=����=���1�rY��lm�Ř�nY�oD����8�V6�u��흕z4V���#U(��7� �,?@.�]x@p^�1�圤?��*�ee�jB�1Ա�l�V��&�H�I��R̷�`)i:�Q�θ���3��ښ�O-a���X�����ix�Wl�d-��;N;:����V�vZ���7A�nۓsvy�X�zԜ�c�N�έ;�^�k���Y<�572Ķ1�F�c��Ms�,"�Q
.֨�;LѦKζ�a�`�sy�a��k@kQm������b7G��1�ڐ'�7����mm��GbYaL�XM6d��[3]���.g[�FW�t1��k;v��^��
�Gm��D�.U������w��<�±����ŧ����`�-������Z�^�҅�gѶ��a�x�k�ZMB�ǿ[��Y��q4��L#��f}��4������J�"~Mƙbg���W��0�m�V�Ҳ��.�iy��R�8s�R�d1'�L����D?i:�pS����r��#j4:�.0�?t�fuCM<hԷ$d�H��H�����!���a��Ү�_լV�g���Z!2�0_N���yҔ;���� "`���n�2�ۉ��yk �h9�alfֆcl���Jd�0DdN�P�\3�#��-xs�3K�t!i�2�N�9�XŅ6�b��/+��تN��>=>�w�Γ��Z���*(���j�DY��W3S��_�n�qwJYb���5A��!m��M����Ox�#��r�U|ڶP���d�-,��p�+9�ޞr�sJ5�ZڭY���-����qWS��O}c/\/�|;��N��}�}ޟ���$�Z�`�O:p�<nK>�t��)����&�0��Z�s�mC
���jIWmÌ+���%i	��B�Ŵ�������fs��ںm������oD�7m�녃>�uI��2���l�����k><;��;Ghe m���a�'�l!2�0M��o�7
�%��dq��6��4��aS���
̉&[�!O�w�ͳ)�H��.1Kų~��#��o2�l����we^�X�"�D�,�_8y�&�S���I9>ϡ�4E,|Y~��-Cƞ1��?q���Ӕ�HһTH m5���q�)M8W[�e"��,�
a�/v՟Cjz\�ӄq����[����Y1�ZBM[5�J�
�V6�4Ut��-�Z�4(�#5k*)�0�ӄe�i�L��Lq���'�ڶX���)�e�-0yM��'�յ�5�ӌ�$.%��8��H��ϙ�̓���Q��:i{�?q�BvR�r � �k�$N�G�q���p����alV{	�5��i�%�F|��x�j+,9!��	)���i�חJۅ�χ�3�-=�\&����>{��ֆ�S{�j�l���D�#��vRd�&a�P�N�l�B[�e#O�|{�8x����~��V7qu�-=�k���|3D�߶��;tg��OQ�+�7�gg�ͮ�;kٺ*���8�йж"8�5*��)A�ґ1��3P��K4�i��*�i��kb��3m�KK4�;�V5K%E
A�$�>�j/�Dx�4�i��*�C˅+Oiy���0�</|��^�lj��C.�<�|ze�VR�K�Ti0��gV3�mCN��oLO�2�΂�
�]�e��Xτ�.ii�3!n�:�`��R��C��l�FR4��{��B6Sq�_#�S���z�}�a�9�
��Z��n��LYOi�
�B�´�aQQ&���*{��*���Km�l8��ģ���jZhe���ֹ���Yy�˫ɻh�[�=����:y�����ܩ��V�Z�S'N{]�k��4��,�M	0�	�.�6�� �M��4�1ÛSX�i�Q�]�[�䤞��g��m�A�q�(���g�n�r[ӣn��S`9���.a-��v^7��\K�\v�hؓ��n�SꃮQ�Ք]V6�6ĺ([�
��~np���ڮrq<��ë+;�t'j�,i��*],-��a�;.�v2J�q��=�'���޳�j�϶�ͱa��
)2�0M�n/�w�zXv=�)�U!t�G8���m��*��SP��3!}�>�fVT�8�!�
��c�B�L��m��ج��o*iif�(��7�����n�#�޷q�i㦜5����A��:C}�e0�2ׄR��zu9�a�K�)���=i�qB�i@�d�ϑ�4��idq��\��F�-�sKOi��]�ޘh��9S�jŊ͗l����cj��H��-*Z���������1�I�1�1���-�b���ʆq~��l$S��=x_��`�u�iB��۲Q��Ճ��y�'���o��N��9��)����۠D�i�lCJ~Ok���1`���dL7k^�Y:�SDā��J''�S���|���x�=�X#�ޖQ��<|m�Z~��AV�����PCIǜp�#���-(w�az*=c����X�q�_��~Uu
G���!
�B��)��g+-�0�u�V���V�ن��xE,�:|����Pi����!)�κ�.4t{sr窞|;�hu\kH3\�u��ֳ1��5��]������Nz|�u��`�i�W�4Xk�t��-<�˛�Y�H������8
e[rA��8Guͫf+����-(�i����Tk S���{A*�0��8�9|��n���ŧ�GY7�Į?(�x�B{�*Sf��q+2��o���H�FJ"P���l��b�#�u�)��Q��B��4�n�����k���|p��S@atbjU��|O>*v\B��`���l�E��r��iһ9S��~�<"DQIFLGR��K�V�v�n
�, g�tn�hFb	D�%kU%f�\�Yv�)1�a:c��}�ro�h�s���O|�߯E��Q-�W�>=%�O�#�Mp���s|���>"��i�����)�OY?=���}ܰϙ��[��E���M�-<�ۛ�I��5�R��P�j�[0�4��R)Dq���.aa����RA�F���+Ba�G�V|��{�˿<O�e�[��Ң��k[�:I�[��CO��/̲�"�R����P��(Z��[(�X����ŦN��a�5�K�L�K1X��1�����3!�3"dnV��/4�����%�q�oc+�t�]��K���y��ϰ��*�8G����#�V����Ӕ��x���AE>P*F8�8�]o��"���)���}�>��a�����T��)�/�c���<t����~�zKU��8w	�-0��sz*=�Usf��H��\�tO�I_��s�u.�2E���sz*4�k˚Z{K˕���l6gɶ�9�O���,ZQ_V�[����&Y�	۷�>'���$1�)MxͿ�1/
p�o�ʭu9��ĸ��mx�l��Yw4�AWX�0����{3�ɶt��Ա���:1q11.���6F�u���q�k�.N�kl�=�N�=`7;��Dn�r2��^�� x���P��Ė'���� *�#���A�Ǌ:��`"����q&n]jW1�Q��:��)�(y�G���;�?������r�tv-���l��bM[��:N@mlڵ�eR-��]����,�ҹj��xc%����p��K��ѵ��3��+!]�bQ�(l[vM��s��[a�	�҄�̛e�,:pqDq�+��p8���y�a�8��L�K���/�h�Ж洑i���w�&>?����ؗ`��v�$�{Lo2m�h��Gp��i���3���=r�Gx��4�k�ß$��MU����.��-=�b�,4�k��҅�V���E� ��f		S��%���8��^q~����E4i��n0�I��dr�4�i��v�U3��;E�G �J�r�y��p\�R�lդ\��>^��W�-kkK�k!V�Ŕ�x����H�-�Ş#O<a��-,���+b��)p��*E(�&sfsl������B�@�-!x=�Ҥ!<`Ţ�ۊeOm��8�<|m�XC��a�L�Q$K)���8��iw �q��/�qXz�عd�Y��_��Y4j0(DL�%E"��~�NR4��6��&{L�y�4VV���P��$h��`hĜ#8�?a�vB8�Kο��F��ڗP��z��[�zW�����CR��Gh�`gZ7F['����������%����Dݼ�3�v� ��3� ����ue:x��״�i�}���V{?7�L�L��{[5�:5.w�����n���p�űI��m�����m;ul�I�=xu�M���Ϗ	�u[Vq�����4���h���G�U�T���p�k���ُ|/5)�+�P�������y,x������%���Ѻ�\;貔	�8Ha=7�8�/@~[�2P_F�c�#�#lK��c�)���ϑk�K���[��<�F�I1};r?�8{��N���}�;50H�*��� l��:G�O۫SC�0���^x�__�����	��ϕ�3�Hek];�����d���	/ި�����y_3F]���g�/Q�㚣~޳Ov���%M���wr�F_�4";���0i(ۻ����NJ�A�9��%��HAqy�w;�AŴ��tȰ��j��鄇�l�ǘ7U/!<Pg�ߘYb��_�������_�����W�u�{Qә>[�佮f߲�'����E�e�9��|Q��
/�L�6Ox�PX��ƃ�{1�����g��_` �L����x���c.�f���L`�?��_?���<��|_ۺv��F73���0��%2H߶f�h�<vE�#E ���I=�c����8eC��0h��q'?���k=4�����X�օ%YKC�+������L"B �Y�ر�d�%Oi�(���qû"Z��sX9���Xk��}�s�6�oU4��{|yj��"V�B��ۆŽ(xｏW�`mA�w�d�7�	�? ��!��f�v]J< ����HĊ':(P��Jō}��e��]�L:s䇽chGȝɥG����L����hЫJ���KMk^M���b�B���~�E���U��O|�jʉ�B
p"��Ŕ�x鸮�?q�-�&��Eb�n��-,��lXz��υ��hj�bdT�|'Ǆ�����Q�Nh4�i��[V�f�0�3�Q?���l��ee4wճ[,X[��-5�B&,��Pn�]�3U�KL�6`��da�2�FV$�q��yN�#=V��My���I��sKI4�}��o�h�_�>���B��18�8E?r�?,�i�w
S=���"��EcqYJ�kZ.�c!� P�n�0���u�)f�(��~�EFɲ�B�ͼ��+8邊�""6�(���(8��l�Ebn���J6�noE"B�R�EtVF�" ������N���_�σ���k����9����U��OMʶ)4�^L�	����Nq��Ҫ#`�-P�rM��Xe�Ō*Ⲫ�fu�;��q.ٚf3�5Xe�R[u4ҳZ�fΉ>�w��:,=G��B,�ź����+7b���8�m�DQ6Č�0$�a��FӉL��)���4_1�&H����8�?av��!& r8�	4�$iF�/�[W�4V}0ڍ,Z{��![�8Dv���u%]%NIi�MT�0�X���E��?k/EG��E��Y�.�jϑ�0�r6�r(�L¤	#4�8�mʳ�g�z�b���}4ڶa����<��|(P@��U45m�Hi�CH,A�~ϳm�.ʵ�|ĵvCj�j�˅c1q-��Fǋ�%6�5ٌ�\�A�"�\�6HYT�[�\z�U,sֻ���7�4.e5t��!�ø�*�V])����vʺٝ�@=�7���[)�!c��c�,�	�.)�Njp�m�5��P-�n&\���Z2źh�E���V�t�a�ۍ'�y#9+;��v���Jf{��_m�Xq��ڈ6��y�T�q����ev�l+�˵��@E�-�fͮ�V�	B���u�mk����F{&ȩUٹ�v�[Z���Ӟ������i�s���&���uF�-=/i��Ti�]�ӄ��r(ȉ����?q�WnŲ��m�-,Za�����}��T�������Kv�@�-ry��Vn�;��ŧ��M^��>�ȅ����Ӝp�gV�8ND���DA:���l��+b��k�T&I��>��}���JY~w�o �E��7�C<pΕBG���є��<eR�J#���g��>���`G�����&-[v�O^�P��ۗ,�χ�/<(E�)^ڕ6%��,!af�ڶ��!>1�H���#�i��X�q���2�#�ハ�t�A����� ��؎M���|��o��E�ʋ�Y�5���wN�!^u�7�~>�_}�+b��}Q�B��0M��o�h��r~""_TN)���r�a�y7*���ݼ�ҍ�+�P����+�B	H�IN�i�O��BZY��u���4Ti��+K����^�����5��S��\U�t�Ǆ�^�/�����K#[��b��3r�)����Ya�!�D�#�ɒ3iGE6���ˡ�����0ښ�<���Zە�@Uvmq�����Ynw�������<���p�+4�YP-=���ql����wfR.�*��:b|xN��a�'Su"d�`�i�W�4Xj7�^�>9������36,�K4�uI���չ�0W�"			ZQ��H��4��S���s��<������/�۪�4�Ie�,�t�ݵ���B�T����QuYH���Į&)�����Q�HaI"p��JTޒh��m�eK>��6Ň���Lb�<t�v�c>��i��B�Zn4��p����#�d8M����M��f��h�m0��9ʷ��W[*��YX勢Uc�ŧ�����O�n��i��דzY��ޞ����yޢڰnF,\P��z���0��=�u��x�=Ѻ�,Z{�n�lXi�.��*b��H*r8D~�zvU���<mSP���k/Eg���$��w��J�1��j$c>g��Õ���8��=���m����k���~ep�YQ-�eXQf�l�a�3L����3\����sC�͆1��b�4͝<'�|��K�a�>�y2�f�'u�_��X����'�?�<a�(���[T\�W5&�+n�d�lAq�����pɚ*�.�I��wP��H˲���'���o��N���[�n�L4_f�&X��u��lXz��][������A�,��=��b�f��ڇPib��T���>)ò?q���$�.2Pf"�8x�
�]{I�F�r��OP�<�L�K�n���^��	���_؈s�:X��ݗJج��nU-=��~�ql��x��L#�<�Z�!",8ҍ$��!���3���<t�꽫>��a�#\Δ-<6�-��,���<�"�P�Komİ� @�O��ު�+�:m�1�W4ƷS�����j�J�MZݳ-�"�5���)ek�K�mU�έ��.�[ʶ�=�ڳ8(N۴��{r��n�*+�3,1 Ф�f��$�ǆ<�#E���Oh�vl�#\��X�m��Yy���V)�˫m�et�f2]Lr��|���w�qkϜ
��f���8�,y�,��`��ݲ�h��{F�s��I��C���-�n�s>X��|�¬��	:�coV_g��\`@nn"b�nT�m�т�5u��lV�f�
DT
8����f����5{J�W��Eg���YJ4�6�d�v���ϡ�4�m2�G�k�-��>5�M����-�yW�/�kNB��E5!�IG=��3���n�ʁif�/����f��5͎�k�I�L@�)8�v��>�m�Ϸ��]�[�W����d_�n&D�|�;�����ggOu�c��ӥC���+��$�-�1�Y���v1�e}�*�:-�ӛ�h���I������ٴ��,���N+��t��c]�s�|�U_k^���Z&�*@�c"B�LD����k>��
<�PA yD��yI><���u��ۭپ�{7����4����Ä��rI�go��\�~�U���U_gF�Uv�)J&T&�*I]*�U};����=�_N�u��Ύ�Qy	I	p��9gN���v���s��5t��n��n���K��8{nj�Z�WB�w2H��+��m��z8��K���aD��`bֲ��`�Ӌ��NR��������rQv���ӣ��F�A�J& �1�yv?t#��׻�.�l���:Qϳ�ѥ����nC A�'gCӕ<�8+vV�~���na˗]�S��9����D�:���˭��݂���R�eA��ggu�Ξ]N�Άܪ��[���o�~m��iHc_���մ��m�X��ܸ��t��]��]���s��zlLyѷ*�y�c[X�M��!���S��-�՛q�,%�/#��}�g��b�OWt��:r�t����N�r�@�AI�iEu����}:�5t����Ӳ��r�ݐ�`L�B@�$�.��vvz��\��h���ӥW;K=ʄ���J|[I�Wc�J�v���8�'u�s�";������P(�"��@(־���~�����eόR(�v��ʻoY��OWt�΍Z)����VH�M��e"TM�MͷM0v�9��3��$r#5Ξk��Ms�f�6��4�b,�+z��ޟ_�w��z:���nU���\P�B!B�
#���v{���������-�i���J�S	( �H�M�ӵ��];_t���z鯣�7����hDRi�I9'ܺ[�>��ʺvw<��gsYU��NJ����B!H�����N�\�=�]��S_i�U5vQ�}X���c���e��D�$41�T6G�D$7���@��!���Y�H�:�{��8�H<�dk�A��]z[����DP�3<P��C)�����l`&����N;3�N��#͟�H�����Ni]����6�tf��O��麪�{
�������</_���$� xz��0B�ZS;[>[v`Ȱg,����F�������'���&����rE����ih�	\
@�$d�y���l�5sy<Om�{��B��K��`~y�.l�zE���	Kh�(漌�1�
a��i��?n`9�w�{�|��=ȋEش�a(f��1K���O�Y4&�!��Ô+���M3���oHsɱ���N4'��Fp���5N�ه�䶴|��bix�1v����؊N��	�;��G�=ߓ��s�5�:�/3���!�-��h§���aƔ)��+g��a^�if���n���<�3x�Z׾����A60)���N�RL�W��żG�ǂ9�=�K�"f>yVW�f|���^˨�{��䇳Ɇv|��161�g=:�����z/<��n����3�Ƿ��d9�u�-gL.B�N�uo�]�C(,�?��\Z��OgM[�6pp9��fzN���n� {��uI�ǽ&4l��8[Κ'h��	����P�q�3Z4	~�Ng�!��eO��{7>pc��UUUUUUUUUUUa��Lnr"q�&wF��wt�B��;n�]��%ڵ�������n�sWa3֮!���2�$���Ʉ���1�6�b��jw �pr`��sЖ����nx-+���(%v��k���>���Ǎ�=��Xx���ɣ&16
8�C�&�ke)�����Ȅg\�R肒�M�eCmF�����a���49�u�Qkb�s:h�[B� d���Ypز�6�Zq��C*]��jҌ��ұM��C6�V�0 �]�p�KZ���K�����2�J[�xb�ݥl���3��l,]-&��^l���pD��δM�u3ҽJ2[������c��ۮ�KU�6<�r�q����.�u� ,-x�s7(��AEt��D0�+nv�c4JĔ+dڙ�C�3b�#����iՄ"�v\�9�Q$۞l^�ĝlK�k R	U""4�b�,��P�'��𘤄h���)e�R˝4�&�V�rq#�7m+�PH0�7�FZ\F���:ܴ�$8�C�n�Nӛ�$T9n�_!�ݸݜ([�<<֨����a��ڝ�mȀW]��,��CʂGMn�3��7)�BXC�G$�I�%�A.vТG���~�0 S��;�$a�^!�Ys�͂<�ft)GX���a���]k4f����;t[���]Z˫�0�v�B*��]]]��Uյ�e�ȶU��b�m4u�Дf��c	�#cZ�ƗJ��:V�V�6�k�1�ʍ,J�QW=
�ێK���a�͜��\#�����'M6���8�/:�ű�vH3smt\�M��G��Vd#YVx��J�m�XN#�3W�#��R�n%�,�`�4�A4tiH<�Y�RG�`��i4m]q�,\�n��͆��T�����9�*|�q�S,m�E择,c`B[L�t�6���XF�ִT�]���J�����f�(u��:��\vJ����'��z������k�\wU�����*�X�k��К(�V�7:�k�>�|�d����Cm0�m�6�]4BjXܻ0P�sr3(��FV-(a���F释�%���+7)�9��(2,�0���(�m� ْ�Zw�j�����c*V�)F�բʅJ�EF���ۮ�U[r$���ۛR�1�cM��}�n�8h���'"�ᬺ���s=N�|�e�h�F8����r�v��y3�<ΛO]�2Wl�ca�LMF���yu�����:��
ˈMk�1ܬ��&�˟ѻ�]��%c[��b�Z7Dl�k-���J�ak4��0�FK�5�,WRk�MX�k��4v��]-���4e� �c��2���	���44*ыf�
C���Yu[b� �D�	4�0e��+Lf�QH���`�M2��l6KE��k4en��9Z&�(�\ed�����?����ӥ�v�<��g���t~�6EP8ڀ��.G"�=:���]uvt�ʪ�j��od��	���ђH+�6u�����_Ov\w;Ou�ӣ�������0c-H��;�J�;zu�,���Wgk���ॿ��a	�+�:q��*�ϲܸ��w]���`#���78RS;W�\�mV�viuV6��1xG��+�v��[3V���ĺ�0�]$�.����gOGԎ��u��tu��m�Zp�$QA	E����oCn:����T�+������#��B�X�+�,�^l};[{��v�;)j�� [����f�Ξ畎�ʭ�+���WgB�h	!#��I}�G.��V�:u����nJ�v�q���@�pE�I���ggs�Oge��Ut����v�VF; ٤�K�L1�M��Δ�Lړ
sL�4���
��K��msj�q�o-�e8�:?t��k^�W��ێ��n�=;:����&I�	��g\�U����u�}��;Hb��&!�@�PF���e����<���4��
-KJ2µ%����a����������M]:P�:�i8�&#$&���k���{���=�+��z��geU��҅0��(RL����Z�v�n*�_�������ӵ�"�`F 쵉����r�����R������B���o>l=�\�S2-���	m��ӳ�%����Ӳ�5�:5�Tl �j�� b�}8Wvs��场>�_N�����ԋ�2I�`i�
1���θE}�۫�N�.v�٫���^$��@�A�a����\�~v���;M\��#P@�%%���{�ngu�RIn1� �{�����E��)2�E")�t�׭��o
�ʺ�_>���}�S�<�hp@74m�]� W�	�6�&fY���Ŷ�.��v��J��J���p� �������0��~�t�~�WN�s��vx.��p����BI#����O>�݊�;:��_g�J;;=iԱ5��)h(rvv^wH����C��uSWgOK(����������H�.������Շ�oZ�Nʭ�ϡ�sTRrD���򖋝��T���:ŵ�?k�u����P ��@��N9<�<����^'�#�}��w�����JЍ�ж9�G73��P�V�\����cs�0�^	��Z���͂����5{��u��G�v��O]ug�/o]��arЍ�2�46���m�y2)�-�j�i�m��Ps�fi��#]�K\ŔL�4�J��~�w�6��e&�O(��(\�3h����!Q�����݅v�W!gm�Dx��Z�ukF�$����8.WẔ��)���`�34�9����l2y)}=�lyۗgL�t�iu#�S��(���4����ɓ:豅̰l(ZL��N&b��1��~֯��ϵ�\b��ϫ�z⸫죰_�D	-	�ۏ�gs�;;=�+��y��ΞV��>�@@��N|�ᳶ��y�w�}�{��z�xl��{HS��Dd��gs�;;<�Ss��p��g�d��i����1����E"����U�y�6t}�N��q�������V�[msO`��&��m��ɢ��;j�ƨ�fXduYkE,�2)ˋb���pXm�y�Z�]=�q�v�d����%��e�Ra"��H�N$C�k�+�����E�ۣ1�
z*�@֩�b�j����|��w}���Ν���z�����QB��Y��s��gvK.v�e�s��坝�{���F?�b@YA8a���S���V�Wk�(���us�}
�)�@�-�"���׆�ή���ݗgo��vvt�qA>D?��M�:��x��<�rq{vfy�[tq��S���vr��R9��q��P�ӮGO.Μ�.���*��}һ;OqWIr�-�i�⯵�]�^X*�m�};=,����à����0���������.t��??����n)nF(!2I���=��J���ς..���.�_���J�!�Ԍ���"T��oNWN�QZ�vr�`���K,�~���I��$��N�\��`�ӧ\��k��zv�h�PAZ~ÅY�`�x2�D��KIyfvy�6x�g��ɺ����x�/�ٙ^y�l[*�:�����������^˄Y��ݜ�z���D#������w%��\���ί<�wb��;O�t��f@Q�B�����gGz����ٳ�NW,�ƌ�Bl%��\����.vw<u���N�;����$��D �w�sr5�����m̈M��K�z�֒ �>��Ȍ� ��c���}Ҿ����}j�_{���;����f�������X�5�쮱8}��_nŝ��8���I�z6�һ�Snp��D�1�]��?d������;�Ys����s��m*�r&��	R����UΕu�_Gm�ϵ���>�+~��H��"���ʭ�ϧ�.>��t�tᳱ����H4\2P)H�t�Yˣ��l���[wN���`���J}-0�};zr��v�쯧a��Y���˝�">g��ĉ���y��7.��%p���HB�����C����Y�71p�͏o6W�H�;����}����q������r�������3����f�l<'nV[n�4��$seYv����j�e<��WT�]�#.&��l��.�	X���Q�6��`,j����[�M5Ы�Ҧ�.��qX�vU+�vf�e ��as6�P����)5��(1�f��Y�jO��h�T��7��������U�e�[�*��w]W&��2�c8vݠͳ`�t�\�X��g^��T�sf�<�X.�4�0e�[�\n���lO]����?��;�?������v�n*�_t��oq8�e,Q8���Rgk�V}�e�;\�����v�6Qd�$pHdm��;oQ���~}H����;o;�ΌwPq��p7#r�����zWӴ�b��ιrW��%��5lJ@[��0##��N�6�=l�;:wb�vv�٪�MMD��#�D@��Ÿ,%<hW�q�\��t��;M21��:.�j��1!!8�S�b��]�����r�ϴ�b~��9�죮����ʌ��y��{׿�I�$�� 	m��<^^�t�
7K�:�]%PD+!Z:����)���z�����`ύ����>Rޕ�T(&A34��U+d�XSw�l�3�ta|*���Zd��9-��1aN��B10P�&�rG��N�n�yH�N�mq�>���[0b�m�B�`��_�?O��湀���?ӧ����L��
+{��C�D�+Z����<:gO��.�⚕4E�V�Ք~���.�y�c����c��ݛ\t��jC�RZ�n�39���	��������`�}�|`��:�lV2�}gŦX�	~����3��G]�Ξ�'����0L�n�����\XυM�al���S� ��QUHDP��&Y���R3�}V���SP(P������x�}�|�����2.!��$nyk�{B$1� �s�`���{���S~�bQѴA���=��e2!��i$=7��ȄQ�YɆ��^!�K�~2�0�#L�zam��[;��M����ob���6ܟq��G��!m���(���쀭❽<��~�64i����4����"|yG�1M����1k���1�{��rb�y��� ��yu�9���p�	)��q��p�3��/f�fG5�0n�ԂZ�LL�X�h��>���,H±����r�'�������� �d��K<��*G��
�t�J�7RY�����SF�E��~S
e�9��A���sb������ǉW�0�RE����9��P&~h�lLi�����ƻ���xc�,�L��L%���AV�(K(n��R_N�AL=0�v\'��Ny�B�}m9�#Xad{��}�a#<_�՛�]c0�	�Ͻ���fk��>�l~��WR��w������O|���t����a[S�����w��g��O-�>��آ�qg� {Wm؇���,��=�n�~���8�W�]e{�~̉�^#"y�=�3c"@AP��)湹�1M�$f�9���q D=Y�H��v�\��>Z�&�=���S��\Ɔ��4u��^���Y��ԜeU��P5���$#����7#��$�DV�Esq�\ҝ�_޻^sp��@�-����E񮳽|`����y�E!6̉�2�����-qc>:���+*u�l�3���T3��~�"J�&�DIUSZ�X���o��o/����ψo�o�gk��-q�0N�\��L��5��ka4�l5RUl�Xf��G6V��c�m���DQyv�.q�n��]A�gwB�yא��>6��_t/�4���ČϡO>����dq��DD� "UI3"f���>;����Tq�ugUZe�9}�_wB��_+��+\tL䨀�QJD�B��_|<��`Ͼ���?�/���-�P��m�M����{)�fT]ve�~<:��q|I��{��Wŉ�7��}о8^�ɯ��&� �wg���ݓE��] �Cyp�wi =""I�ߪ����W���W�.�%zTUN~0�,W�|^Bf���I���숴���,}����]��#M�ËD��J�0tc[���e`���`U,hJh�R˯6aCh��͕T��Ҫ�����ϊo�U���T�t+L��d'C������:Ϋ�*0��"2�D��DUAS35U7�Ë��V�C0\���|Y��}�f	��ܯ�iwL�\���f��S3Qk��B���/�8Xu�wE��>;��|)8��>��(g��}�Ԣ��UQSH�0D�_>����ɾ0L�z��}о8��w´��Bx㾋���r�ꈩP��R8P�)R�
|U����0�8k�a6���	�Gt_>��W}8_&���@)��%IOw.#h��{�D $	� Hp�,�� ��������lQh�[���۱�l.m9�n�֙���+nQ�
΃۬���9�����h��v�Wg�����뮉n��ť��k��)
]n�cH�m�D�Lx��ڗJA�f�ekn��D�Ital��Qkv:!*�n@�����ܱ�Ӥ�È+c�;f�%䵢�jv������Z�<v檉X5]5�hk�g�:�n��m�y�]oYtSe(LU՘�`�ʸ�%�\�pv�7oT���LX^g�m\m�e�-���8���[q+.rCV@����U&�UQS��������Ze����;���������y	�<:�o�'�9�,-X�մVN��?��ǿ���>��}]�l�3�+{�o�Y��u�qk�i�B�����'�ILD�nA��?����V��L�_nM���|��>#��-9����D���!(��Ϝm%5
�"g�>��}
�4���m2�_Ц��_p����_P�����*��!5Jj""f��Y���-2�|-��W��i�d�,LÝgz��a����G0�IEx�1˵5نՌƴǤ���K���9.��re��&����ΞI���ꘊ�-3gО>�����>��e�&|vWq|)8vL�e��U�t�H����L�""*�Wŏ�a2�|y�^��@29�u�W:tۛ�f�+��{��c�%st%�TZأR�s���S�?��L���&�Ϋ��O.��R���S4��e5*���ύ������m�(���\�����_�y6�>#�\�-���آ�{N{)��k�͖�#/!5����8_����.0���_0���ꉢ�b�1"���V��0\��c�X>�2U�ύ����T����Bt�P�cbb
���s��_����<-5���*�v�"�d��um{{C)n;:V�\�g��|N������&�3����Vq��운��o�_wB�y�2E�H���*bj��0}�?�a}��Zd�ϡ<yԯ�8_븾'!3�_�Ȕ(��T�(S3Q|*8��ݓ6�c>Ow�����X�)dRB��r2&�GNgw\�wt��Pc"s��5��(��L�ܜ/��t�t[�Tq�1V�� �~R5�:i�!۟��Ƽ��y	�����⶟"�3�F�OE*B��IS5Q|P����&قf��6�i�yԭ2F^Bk}WŜ/�b)wTz������
�f.����
�Tl�m�P�\�x�a��lb��F��ٹQ�V�1s���Bg�vU���z���f�wu���gt,U���&|E%GE(�����&j��B��.��Čϡ_>��(�|t��M��0��t��Iŝ)�(�*S33%*��������[7ܯ�;�|Gu�7ŉ�k���}�+����(e�
{ܣ�h���$�A蚚/�8_}��d&|7]�|,8���k��ăJ|p�H(���[����:O9F�9IPRQ����^}y��u��l��A$M	MU*�bf{���g>��\`Ͼ�u���'�E���gON�r��70#6�3ͦYY�h�bB��ۮz3�R��>Mn�� �8�-f����fHT�T+�a���>E�0g��}��Gt/�}E�����o�iV
�Ҫ��P������0g�	я�������&���ύ���ËW|�OǇOH���pQ��m�y�ú�2��ϊ}
�4�}��P���w�|Q���F(B:�b���TLЭ�p��7�q|+8ú��\X�y�W�дu����)N�8U3TL���"b��_t,8û����`�����|Y�����]Bgŷ}7³�����˕%w\�$�K�K��!�Qb��9�˻��L�9rr�i	�HHp>������k.F[8{�Pl.6�g-��n�7��\e���j�w-� �r6�������L]�1��dҺ86�d�em]&W��Me�x�]�tqkr��vT�i�L��gո�m��9��@�f6��c��]����\��D�*�I`��L���#� ���n�v���a2ݬ���$I�,ntҶ��j��]â�:�Cax�l��l�D����I��l�Jۚ����������VR�v�]����o�u��'��m�����M^�յT��`�������-:s���!�t�t*8û>ʵ���W�]�Q�b�f �"��'�X�~��_���㾅|,8�����������N�_���#-A�ۋ)�S⨿���,8}��qc3�N����g=��T&ao��Tҥ2UQ���5�Ë5�r�\`��/����î��قe�o�/��C�&>��!ME)��"j-2�_Э��o�8_o�e�&|v>X_
�0s��6�C0U��� �Q��ş�n�-�1k��U���{h$�k.�j�Z������n7;�����0����e[0L��\[�Tq��.>-3_Л�;�0�|B�;�SQ�L���$D�l��ϋ�}�V �x�:�a��D�db�����%�\�I@n�cd� >+�dŮ,g¦�0�,}I����Bf�r%�j"bh�!J�B��;��\`������Å��Y<_�������Xqdo.�J�B����DD�EMk���a|P����-�&|Wwd+�gWwх�X���o�%}%L�")R�57Ŝ,#�:o��L�5����͛�\`�}��|a������D/�R������!G�T�efv�	G
Eu	��rZR�#��;YsR���l�'��I����������>�\`��]��E�G��d�&a�r;�L�&���&j�_
N,���L��-��W��i��e[,LßY�o�a����T�f"
�bQQ3E�X�����|Y���]Ų�k�Q{�r�C	wt���
��̚H�.]6,@Rn�TX��
Ȭ��1���7�9������c0\�쪅
UDMT��*��_wB�{:0�(L�;���B��}�M�0f}	�>��:�b$8!U
bb������*>/������E�Xυ�]��'t/��M�ύ����A/4�8�n�<��m'=�mgny��9�Ar\�U�Le4�˯V�EǈR$��LTQ}Ь������3>��?���8Xwge_p���ɾ|S�_"�zQQ$LIUUi�3�ow�
���/��^J�`��]��o�QƑݞx)�NjM�<�j6�q�YQ8s�㯺p�]�g�7�q|+8��gUZ�`���$��r�}^��"JAJb�D��&a����0y�|Zf���}�l�<q�|Ut��AE�w\o���̪$LQ����2Z0(h�M��J+��LDC	q( ���&�3��ɞE*���SRELUM���{��3�>迢���,'����bf��6��|S��ɹp++�n&��}��sMt�� Z�3̤m��؉��5ΥA3E��uUD�U6��>�;���g
���fd&|^��W³����\`υ�`qQ3JiMD ����X[���bg�S}
�B�������3�>/�o�8c�Eg�ѤZ�@SeI&S�
t������ou�3i�3�Y޾0뿥[0L�)��#�IRI0J"h��_iwO��$f}
o���N}Ӆ�w	�����:�/��&�h������3�.i�>��%}�U���;�)�V2���B���2������j�����j�����յ�U`��!�h� ��Z�_��տ��Vm�M��UiZ��ڛUeki�Vm�J�fմګ-[M��mT�Vkm��YUi�VV֛UemiZ�֭6��m��VVڕ��mi�VmmM��mT�Vj�mU��ͪ�UR�YZ��VV�6�ͪ��ejͪ�ڳj�մګ5�����M��֦�Yj�j�UM��kSj����Ym��YZͪ�j��e��Uf֛Uf�J�f�mU��ګ6��V[ej��6�ͶmU�R�Y��Uf��VmJ�e�ګ6ͪ�m+U��j�՛UeYZ�֛Uef�Y�mU�J�e��Vm�UeR�Y�mU�ͪ��j�lګ6�Ue��YVmU�M��YZ���Ue�j��6���mi[mkj[m��f�YV�j����VmVmU��ͪ��lګ+U+U�j�Uf��ګ6եj��u[Z�_�j�� ��� @$! ,B�B�$! ?�B�$! ?��!�H��B�� �����)��csX�Ĺ,�������_��� @ p��  �J�   Q@ (�"�I �C@ �T
]Ѽ > �� �@�) " JU @��
  �%�Pww({�ض���
B�:{��������h����W�W� �ί���蠳v�t	c�]���֔�E	}�@|�@=���U�mI���b�7{�ZS�UW@p	҅2ݫ"'b���pS�SN����h ��:RK�� �*�l(¤Sʩ�J#Z��u��j��v���v�^���5��^�plR!li�Q�P�r�&��v��@iU=�S�Tk[,���Y5��ҽJJ(�X�B�K�.F�At�(q�`4A��5��JK��U�[(�R��h�j�=/s֍jUvl9�9���*��W�UH*@+l��Z2t�;��V۳U�PH`=�W�����o3:eW6��Z�*=�C�����	�)J)�*�="��M�R�`
��d�����w�Y��=j��ws�*=n�*�P��T��J�PI�t	��Z1�W��OwuUF�C'��0�MUw3�z*���z�E4:uT��� T�VrG6����TZq\�y�n�=��q�Iswj���w �iQQ�1�( (b�uր;�����J�2&�9
֨$�J���H��W����Z�4���X�V�(�z�r*�h�hj�Y)�ѡ��[�U�w@+fQG�v=dS�                ��T�S�4�      S�a%*�6PCCF`�d�d`L&���U!�&��a0�L шɈ�O"�
���ѣM4ɣ�dh4ad�hd����@�4h ��b ��$�B`� M4	0lS&�"<�������ͼB����k�cEk�7�Z��!���8���M�ڊ v����E�s��ae�eQ󂢂�������h�%�J"C���ʊ���> \��������_����8�?�В�����C<��xX��h��(X�\Y]V�S��>/�t�ˉ���]��k�re�"	���x۰ד��_}l�!�q[�"wr��t�)��z��@����Q�\�]��<�qJ���b��e��t'2#�x��A�ʜ��ӠU�os��8 ��$T�F"���1�<�[9P��$�ҬJ�= \c �㬰C'2���8��H��U*�"q"� !�pK@�S�)P]D���2���c�	�׹�_�q����q=�u���u���/m��$q���6�w����l��~���_�~��-�{�Qs5 DC�Ui��=�����y��	L��z4a-��m��&�Zzh���ԥ�A�Ut��*ŉT�����/�}G��>���<;�	�;�ُ\כUz<%����`N>�P����,|���5����Ж/"��~b�p���#Zu#72�v��) �7K�i�[���R�)Q(�ƭ���_n5��?��za�!��(b��^��uل)�<�8a�6��۝&�*�	8�ٽz�Z@�{����-�Mr�c��Hz;��ٿN�N��G��i���o;d��Gi�m���3��KB�X3� �+ׁr:��ĳ��ٶ��
��XtFܬ�{4ޅ���c�^1���wCւ�GBmCama��y�4��$�aP�;ذ�3$��	R�`9�C3PTƉa"���g��yv��5Qpr��kd�hb��d�s0Ĩxgq0%�8D{�{Շ^���b��N� Ӽ�qu�7�0��ۑiE�#�ې�t��EM���׹(b�V�wC��˪j�B́]\3QZ�I �<���Y��.w&��
w���PU��T�߷���7Ca�Ef�4�U�i�K��Ǭ����Tw�C����i��"o��Ig �7d=Yx8n$��3>y5ǲ�������i
[�w	ך�*�����>���N*�E�s�A�������=x�$s8*�~�JPJ,���%k���ָc';�8��� ӻ��š���3��6�o[���2}�&���������N�x퓶,��5rzާ�z�c��1���e��{���g�Y�v��d @Ƶ�����v!lzoS�{�yVk��eSTX�h�)��r��<�L���gR�h@4Gѐ֎����Dj-ہ��oV�J�qn�P�fǗ�#z���y���euv��R42h5p��Ov��������	b��c9�1Ib���a��͙x^I��l^�6V�];r�8�onv:��V�e�~9�f9�^}��v�����Oh��.'+x���e<�Z
(���wc���{`@�XICXc���x�p��eYӇA��[^>�g�vQug�,��0��sy�S'�-]��C���p�"���ɖ͡U)Ʋ�v�6�Y�1�O�/��y|��4MN�7&m�<��':[����$XF�J)���u�ݬ�>���w��M�|������#���X��6u�s��H�ĉ�Z�*��8�S7��xr����9L�Ȩ�c�Ĵ&*EKD���E���'_eh}fv\��V�a��0����^iãuG{H,�u�6�Xp���?^��ر� �@���&�wH�{t�/���g$�׺Q"��hR7�;��~p�up�sg��b縱v�<wG6��:C�:v�p�۷I�R����t��ɹx8 �'�:ɢ��׬�;1�|�{�r�#^�T���wh�N�vi`��WH�wH�Gaj`�|F���8�W{=�^q\
ocUVC��[��g:\p�8��:���u=�M�&�~��Ӥi�erس��z	�qC�R!�w�P�n<�$�c�ˮ�R 6K���c#;0]�MZ��n
�,�Ӈ�b�ئ��^��\�X���v#7_ f0m��S0���3��5s����\0�u�5�W���!��ĪiUҢ���<2^��-Ʉ��r�~bdg��b��w[w[N�!�^�L�P�#r�q���xv��.mb%���	{��D�2Pu�{�ѝP=5�91�9]B��$�;�kB�i��U��K^(ʽ�퍹	���[�V\�� -f�B������9�U3F�ssr0��Z-O��!��,R���]�Zz6d3�v�Ğw'5�3d��L�d���ey�0�+��m��K�q����c�Ȟ��e;o.��r���dY�T�l�r�:w[�6�}��D]{��4�q+9����%n�tXxw��OAy���W/����@�׬���xUA�;fԦڕ�6<���8�������jn>)ח��-�Q�D�pǈ��F%�N��A�R�M̧��bT��+}����`��N���ݡH���B�˺P|�͎�ԛˠ�i}Op�|l�g:���n��/�e72� "��E�ݻOot�݅�e�Cdm����7׏��hTC�(V����L��.�'�����%U�j��l��6�*6Xrƈ�]cŜ�@��%!ύ�.�uv��w�^�,��QbnB�Ǯ�� ݡ��-	�==����gD��T�N���4�w�Mf��Vˈ[�����iu��Ռ�&��٫6�aB�eѩ�d�&ʹ�fjت�nx�hm�"�vtX�������gGz�*r�p	Kq��]J�ߝ���4��4��7U�Tm����+��$��W����s�FQ�A�U����z�4��=82=�c˧%�MYM[83Z�&C{��J+*ȹ��L1�QwV�VR��h��\e���rs������]��y�sT��Q�Vs�Yχ2o�$*�p�\� ��Z���ԯ]۴�ea��pL�y���-tș��D���ֱ�ol�3�n>�\sr`(&�q��ӄլN�g[ܽ��/N�@ͨʹ��*��L��Zy;=�ϲ6[�(�W��My�Ns�����r�1@f�"��I��z��Զ���I��Vr�� u���y���!�ȍ<�E�%7��sJYt-Tv2��s�yy"���!��;�-xӷ#��W�<�(�坚�gIx�O_Тa���n��[�L	tv��$3C������ƽ���v�d�Pyc��ut ;,M���5�Ob|��i�[��q{8�ǭð��ż{����C[ř���T�ܷ��֒@I��D�R.ذ7��:�b���,+b�:�3���7�i����X2�Ӂ.:��A��5�s�K�e����wJ�!�&j��ƚ�A�*{@�_�՜��t�Kr�ͮb�6��r�v�ܱn��;(�R�����p��8n���K���y�J�&I��w������3%��Z�+���f鋻VC���dc6�®�ف��X�HD�|;�=�x˸��X�A�A�Wf@JnL��R���pF���u�F�+yb�駸���F��9j���;6HF�mWeK�w���0yp�F�8���*;�^hC��T�ӥ,ۇ�8����7RSGa�m��`mr����:���ں�;v��\�>�w(��z����T㯴��b t��LۯN�82?3�ݑ��`W,%Dn��Ʈ�k�����C#�����F�I�.Xte�Y�۸��)�]����CQܢl�6Tӫb����E��Ħ��;hޒ�KS��@nkȑ�glzs]ǢZf��K7)-�$:�U���s�{n��y�nՍ2�n�-�te��ح�u4�)E����f��	u�^�Obks�J�j�8�8���#9�c�G6�&�kٵ�4�o[w5�;�aX�Ǐx�Y�*��I�Kݨ�RM|+�ͻ�qq��Y>A(��Au��<1���X]��f�/l�\\zcn<���������e�R1��')���P��os{wA�ǽg?�]���c���9S���n��`���C*��50�}ڇ�Î��=oV�21)��(�/]#��.�j�k-n�n=��j�T��:���kCh���`��qLU���Ϧ�\xjVǵ�ɠ[�k8�"�W:�N��]�ZY#Rq�\;���Ӭ�Gri�Q]�۫�6�!�9����S��T7��π������U���ڝ��B�vQ����*�6C�~�?�p�6sn����f��?]d����?7V!	�:���I�����`����U;<��\<�j��E�\�<m�u�3a��)�X�dF�r!�:,h��g� �H���FX�4pԿ�%�T                                                    �                    /������|�������GJ�D�D�T�mζƖ�ܹ�ū��`4���m����hvB�$�P��q͂^i���h����JF��//Hq���]d�c��{�J��kcv�pK-l������B���t�V�v�M&ˬ�ee��mq��UZ\@䭊S"�	���S�bX�lt`KB	��[��p.������_��5vo):R@Z�.��.0�)Y�]�s.V&܎��$�u�Bjsz���k[i6V��7I�e��Z�u5��g�qo3:e�i�֥�N�f�/Y,0�vh:�/���omۉ��#R��CP*.٥��App���0W^u�.G$��ɰ��u�u˩;\E���b�0�K-�6�!��gJh�ma�1��BĴ�]5lF䥚��Ҭ������ml�k6;Jض�ء�m���$��el�^Խ�k6v+��#�9m�cw9��֪�����b&v���X��� W2�]��If�cS���dln+��1�v#.�%(�����Ij�_	��_��%�X��)���F���ems�nu��WZ�ġk!���L����x�jV���
dtv�ݦ�Uή��+�7ku��x�"֥!Z�l��4���Q�)JgY��`��q�Ie�Y3t�)j�\7],���A�^k=&��f����/r��R�����zݲ�PfXY��;\���k.V��5#)�0��h]�CD�e�R5�*	������cf�Y�eBj�H�Īc �/`��.-M�r��6�r[Z-԰���b9(��li@R��;]a4�Bt�P�X�v��6��Y�,Y�PZA�]dHlLnڠ�6�"C;V魶����J�L�f��Ŷ��w�H�R��ӷ�
x��D�6۷N-��\uڮ;)SFi�::k=7bM�n�7fۆnW;�p�˝Ji��� Z��&�q���&j�VԼ�F�^۬��L�9oY��il]J:X6b�A�,���cD)fj��-i�.��XR��
�Z�s�e��֦Z�ä��YMy�����ޛ��F�/[��k'����-��Z�b�dՍ�[s���f�1��)j*hFT��Z.r��i�X���Ħ��SMر�ك4�:�5lٷZ��iD ��]��E�6�	���F��Ȑօ��e�F�ee� ��YVŮkG��\�]%m�Ĕ�*�-��ݫ�T���$��[6cvͱ�ck޶7�Mt�Yp��%";]u�i*J�m�;�1��e��.c|/T7]�j�w7m�lnvʞ��ݴ����Ӧ�s�μםUu�kI؋��&�n������W��W$�ɴ��u��W�JB�-�2���5�	/��uۈAi`�j�Yph�e,���ٰ�m#-��Ԏ�Բ�hT���i]
]3q!F��:¹�0iV�!�c�n�	ll�����؁JVk�l�5%�V��`J ۭ�x�R��ƨ�6�b����К���&��K2x�	�|m�u�&
ٵ.���f���,%|ω5�VSf�V��	�y�Lv��p9K
�7�ЃE��6�f,��n�hn�J��$Vd���Jn�Kd;7t弜�7&�gG�eN7k/k�_g+eڸ+�Fi-���Li�F��:�h�#���m�[m7٧^e��1��}�f��dN������:�|����ۡ���%MCn]l҆��
u��Z�vT�v�:�gYEf����J8)����b��.m�yz۩6��$1j�۵Cv�%�F5�ݬE"V�mil,Bᣇ'f��h7MR]n���˫��q1��:��h	�Jj+6ڔRˬyu�.����X�̥֮�� 4x���(0�c[�Z����r�
�ѩ�T�0�r�Rj���2�D�U�ۊF��MSWL�4�Dv�Z��%���-٘*�b�@e��R�anM��E�F��V�#5�9S�wgb�vZ�@�5-�\�.��FLw���'��R�j�M�u;,6�\��Ra��u �.Yf#^�t�s]M�=gU�H������,&Ј��ŷ!M�����+Bh��3-+�&�Ԛ�0�8�hց���©�h�5\1�*�i^6���]�M�6ʁCZ)UP�Z�]�ƈ�m���qb����K���95�:	I�d�YG[��]ka4ѩ�L�䅲��ˠR���9��ignz�h3�.Ӥkf�m�a6[cEKt�e��t��]�Yn[Z��ڊ��A�d���ɧe�]{:��؛coH����a��1��Ŧ��-4�&���Mn���̺d	��dI�YK܎�;�k�첅�]�&���3n�`�Ͱ���;K*�k3��T��9�	�a�4�X�dE���&�;m�n��i��<�2�	Wuk(ŷ�g@�S�N�/�/,�&�\q{NҐsnah
A�nSm#3�b�..��As��iI�iYj�e���d3�l�nd�[��+[թ�*�Ɩն��B2���c[�wzkUf�o��\�P6�eP%���	�#f��+5��\jh�̰�l֗Ie�ƭ��Q�&�&̽v�5��Y��]E�]�n�"��Kѭ��MY�-U�f��&-cb��W�A�[\�H�Q�RЦݦ��f��eƅ��V5h�okbT����!�՛/Y�l� ���ݠ]�lc�
�����0���+aX֒�����Ƣ,�$�n��m�\�#�]͙�X�B��!\%Kmm�P�mq�ju�d%w֕�d�"�B�+Wg��ZR�$��x�����M���:;X�j֔&���^xƅ�F�4�Afc:\�k:��y	�[lǵ�u��&�cb\�hE���ft��K ���Zg2��m\9��4J�#�&����Y�Y���s
����n-h��5Y	?��������w������f�#���wj���/�;#��<{�Z�z-��|�ےIsik�'�PUP0`�W@}Q(ɴ�X��Kڎ"`��=rqӫ�  �s�^���nOy�&Ǜ�
A|���բא��ܹa��> v��%����h����~����@ D`���2z�]�u����@
���|����� "1"I?��𺹏�-�B`�%qT(z�Tgk��%q3��h����X��P���};����|�         �   K�����HKk-�,�
J��f��aMp�X���R5)�L��g��L-�f�m+UԖjmc5T����钔�v��G��,�mc5ڵ���Y��(�f�Ү�0X��Aչ)3�i�)L�vt!1P&H��4�M5#�``��.0�o;^E�Y��*T���o[�'t��1,�^�b��it�	Z�rP�֪LAC�eK�Ɨh�6���3�n�f]�����q;v�`�5a�f5&s��h�6��#5�@�&�tZm�<���\;��L�
ኣHQ%�kRY�2l�A��+j��{�l�`���%���ݴs]��0^Z�6ljv��ms��ײ=3��u��%��5�9�t�Y�a�c�a
�T.L���vb�l�v�;u�E�S�]���n�m��M�nds��7mlN���m�*�%nk[14�[�툈gR�\8��q���7o^M//��d���mr��Mjb�	������XF�-Mm�bQWd�Jb��콭.��k����h�k�/@��V4���ݬц����0:V��$)��7;MG�M���P����������K����/�'���̛ܱ30^�P��X�7����K�? sMz�Nݻn��͵�k,�a�4�T5V�e��WJl��R���دdr�m�՚�ic�_Ix�7Y�2"U�ʸ��B�qBfS�(M��[�#]l�{9yv�H��+�ԅ�,�6y���<�}U��������ecN5�%-QU����>'�	q{�"iߑW�A�U��ô^�L����5T~��P���n�5��s�)R�x��7�M|�>~��.����0[��z�n�#3$�!:Ns�d*Y�Dׇ����Ǐ�V���b^}p��a�vt�k.?J�X���3$1����h��T(�0�e_�R<j���}�`�X��lor�^�M�I��HʅJ~�C�fH��!sw����j�l�Eo1�:���㈳��&H^���Ŝ��bB��X�s���>s{n_���eF���� �Y`��Y�Z.?�E(�NAG{e�� ��N���b&���:��&��,�,��ӄ}��T�z�~�������Y��v��t�,����_�Τ6�(+�F��\���!�ʯj!=��j܋�̬_�~h���G�GTk�H����6坹��G͛����풯;���=��~����]�}�~��������ys����Z%�f$UF+�0��`�& ���l�8��m��-����GN9|\�K5�3�8�A-�Cb9�oT�`b9��_P3���x�"�,�mF%�g�j�P��k�Yd����$RA/A�{K����M�M\�qX���d�UF�Eŧ'_Ȓ���X�L���. L߂�gjoC1d�(@��*;�a/Z�+�w�m^�b�}N Z	 �xⱖ�ַޔ�w��"���[����X�>�W!�� ZÜ��P�H֕��3�Z�N8̈́*%@�1�������q���uPoQ�x�)���/`Kʌ�TMAm$	��%��H@/������Z��7�_Wǐ�Y\�b�nX���@+e�ãJ�h'u����V|�|;��I��LZ������N5,x;�
��h��[m,�$��ꩱ	�CQ/�ٖV�ێ8Ε8���Kқ��8����q�c	�5��8 'Lw'�:I�~G��W�6���3Ih�� �J��  "#������4���?�� �)�/eu�dF�v����B�7�X�MG7����x�B�qi���ILml�X�5j	h�@���N�#N;K��%��q�]����fb��w�|P�$B��%�HH�Ƹ�!�,�3 �KF�3kp�x�K���X#�_�t��"�ٌ�R*�]&̪;�Jͬ)��r���(��- �[@�9��4��:�
bU&f���w�D����Gx$�Z+���[mz*�X��[(���V3��zα�b�q 13�m~/�%�5�dWk��h���$o�W���T*(TK�ͨL�"��V��4(o j!���/�v��K캃x֠7���Z^m�hf _�8�*b�5�12Xq.ƒӋ�
b��@L�{U�@�2I��IjE�;bM�3����3D�o�giH;�R�[jY�#�� � �Sxc��|A����j�x�A6���6S�I�q�٬pJ/�in��2�(���ĸ�Du��w��Y�OҰ�ޝ��q)F�I1E��8�� �Z��EW��]�ckb�	xg�x!�G7�^#����UJ��`��҄�&aQ���!V�Î1k�� m��D�h;U.b�C[�(�t^I�F�	�P�P�Dd@�*&�n^�x�#�	}M�kkY�fP��T�fY	0ul�I�jJ�b���Ve��R�(�T��(j q�KA���P�_8�K���X$�Ix拌\W�_G��N��0� �	"6��q���m�8�f��mN�����*�xb��GQ5���3k�0��C�zR�Ә$��R�
.'=8�9�����J�zA�� fZ(H�������ե走���L�-�jZ��|�mD$�^6��r�Z��^�A�$b�_b���֩mE��!�]�f�X35M�!x�{��ۺU�^���2�$�����P�N��;m��esٻ�ISn���"��p�4����q�[�qO�ĐR	=�{�O�6��.1s�E���qX�m�W9���W���u̪��^��@gmd��5���Zj	�LA�P�9�7�����5G9�x�\��{_w]�b)	�NT�)��f��]�Um]�iH�B�f�%�k��\g,I1Q�T.HZ��ad7�P�:��/Gx^���涊�� b5$��CPw��x�lfVp;����1^1X��T��c9��7�b��$��XN q�0W�������)��%[V�T8��B��I-ϵ�y�I(a��G	�!�8�Ut�/-�o�����}m��b�G0u�T�~(�0	z�[qm��A8�I7�7�K"{�Z:�t��H�ΐ<9�����s���^!Pw�ʍGx���a�0-��X�UD��%@���B��i`֥%����%gk���}�"�!��!ќ	���k�؁�o�Tw��d�q��^#P	�/t$K�7֥��L�*x��/�8ߍV09*�j�/eu}>���ėo���u�9�֮>qx�*0�h�}��h��#�9�H|s��@�x�Ƙ��	>�./6"�s�����+�];���Ӧ��q8�,��\^�B�ObU�bÛMq+@p,�=^q/	 ���P��g6��~��OZ��.��g�ʪ�+[&<I�9��oep���S3�9��I$�H���7�{ӯgN���괖j��k�定mt�G�hJ�%�����盙C̚[��p��65��tܰ���3�]Z�-�$�4V���i�	��KrJ��є�l��S8]����6�tz�\�Y0�k�����Ѧ��䩉fv�*���?�K�$��Ժ�r���jD+j^ ^�����Na�v�ŧҮ�=:D��Vwl�ll���o�	���F��b�{Z�oY�8��ƹ����i�Td�1sNAs��#q}���� �����&�
���Bĭ_��9��/�sE-�|C���Ϟ�A�0�S���>*��招��y��g$���(��M�!|�ӟF����	/�&.A-���K~����E;��Ň���9e	@=�%��{�r�q|y�Z��4I�Ę��%�t�Nȴ拐L�8u.���s��|��A�����s�߾���Kk%
����|]9��b��:r�ײNh�8��s�Vqz�&+,�b��\�,��t�mL\������B�P�~��J���_:#拨�[ �R� Z/��Qģw߻y�.��Շ�NtAŢx�-�-:(􈨛@������}���رx�fk4�y�t���/����u��n��]C �֦�ZZ������B�ټ��]���(�7_�xX@E�;讟(����NB�+_++����T������e��ӧ��b_}@��T�ۿk�0W����	g[�8��_yOr���Z����]�v3{���R�o4|A%�'v?վ�Z&x/q�_�E���KΧ�g8{�`l��4����>��?
�7ϖ�Ծ���Ӑ�,�����|i��
��/�	��a�@g��K�,Q27�����~�9�����fi�Fő=��^���DB��҉��b݀�s�Tz!X}tF����稸EPqD����"�LkH(�|��V�9�A]�U�׆a���+�ou�WZI�	��uʔo�h�޷��ǚ2���Σ���jӽ�~�ig�p��Ŭ#r�>x]����\�k�D�M��(��(-��f6%���>+R���x��Y��-_��M\}t֐�h�LK�^P�6)E�=չc�e<\4���D�`>���>�/�/9Cx���!f�475���[xdI����[~4��������zm�0�<(������绮��M��3��:�o-�'�ժ����V>m];���An
��Ֆ�X�C=��<��!}���1d��u��[���w�trM�����mhȭ�w�go�?PЗz�h<�����y4LIf�va��Y��:�;,r_g�S+�|�h���5����gf�i�|r�mآ���!^𷰹�+$��M��c���0�U9�S�9^R� �6�G�R|�矁��	���W,��-t
1��Y��Z�e�S�	[�#����o���YB�"�[$pS���=77j���g�-���'/����Hd��Vc���z���(�7��YY�[Ĥ��z�:�_-�¿��5�G~�*)I�0���,JY�pҵ�W���A��#�y3K0�֫�8����O�X�jb�5���y(ME߰�&!��E&��+'���q����"K�L�߫z/�����;h��nˑ��+��ޝ���.�[�́u��IB{�g�#K��+|������O?*�p�5~1��e�9ش�$aE��}&x�}ތ����.��7�3v����\|��,�yP�?`?1����i�K���<�qf�h���l8�d%�*�~��׬Qyn.�K��ye��G�]�^�Ra���rn��p�H���"F��D<��E���=�g�l�g ��k�o�����f�b�a~��Da�����|�>�( .8i94ƴz�x�G㹌��`�����gf�A�����?�Ӫ���(b%JA���P�h�z�}l�� ۧ�&\�u����8`��B�"m��<�S�$�F�ӏ��[��؉M#�L��r��k����,����^�r��~��}t>�0{�~��'\k�	����#�:{��Â���wJ�ن����VI$�I q9  �i4�[-�&
]%mfc����rZْ��.��W#�]aL&�۰6 j���Yה�+�ky�Ss��T�@i��Pډ�,��J3K�+�ζ�h�)�
m��5�u�+Sy��ì0[��bEe�w$]{fU�"�}�JR)�0�z?���EN2:�w�ˌ����z+?G��d�8��l{dI��h��M䲯i�x�-v_�w�m-��5^�����j�TMʶ�ƚ���������N%:Nq;ڗz6лdkguMB�����G�����R�0����p7F�&a)w�G��L�m-��1���x	�;γf1.����񷏱mk촖/6#!u��s���>ys:����������7���6�l�$� ��u�_����E�n�b�h��t�w:��D%�فA#Q&s�0��5f�]v�&j����q_�_5�,�@ƮП��no3j}��F���z���r��dk�w��E��r.=JʮT�D7,X�Y�.�΢:�me>v����Q�-�r�|���~D2�9\�{�l��/A�O&8Tl�29�l܍�����vc�����C�����|_NI��O�2'�T����̟kP�E:Kz�P��M˒;PTA�m�B�0�7ӶJCsr�o_n��|B�~�k����&�;���D�{���3`K��գ��d����㈶
��[
���Pإ������f�-�|�Mde'����T�=6�E(��7�G�&XG[ӧ��rL+��� F���L\�p5dՌ,�N�9܅ֺ��ᇶ�_5v:�J��P;B1(ɖA�kNYXF�&Bx��̉	ZS����/��n�CO���,�<�� ��H��/�*�9��^&��k�nW���k�j���fh��;�|3M���C�}��������+�#�¢*���'�YvLۭ��^źgש�nG�_o���C��� ��¨ts�*����r4��B=���0��ח�Txj��7�����ҧ�$��SJ�nv/�C�=�3��Hc|��I��$i�=���EsVļ��yy9�K�b�3r�9ⰻ����$�쉲�udq]�X6�ヮe����[/p��o^,;����S��G����B�w�;T�q�sW%h���ֹ��D3װ�v���&���GC�V(6�Q��ɦkS]+��_+���yk�l�Z������`��ь�Gt_.u��sToe���Is`x�E�W(���۾<�tўx��w��G	SZ�$�W�7����*g�B��2��Ej͒�5H���?}���׃��!��#�'�u�n�_C���%�����0����n��`�Q����׳��G����2�q��]�)��a� X=�i
B�}S��>��#F�|�� .B��[��\e�J�%'Z)�";{)�v@�Y�b���?GNt���YK���{R6�a�$q DH)�z
K�]s���H��$�|�;Z�N�A��ˊ�H�<n�Pw���_�;Z1+A�	 ���f�N'����"d�Lu�Y��hᱎɲT�\F%|��^5�C��y����ٛ ��9;��D�?��R�I��	ì��Sf�c�wy�}��}���wT�]W!^���"�ߊ�K��̶�XBmէ4ȏT,"!F5�Z.�KD�l��N9-Ύ�W^�"�fù��m[/E�5�p���$q�̲�y���zx���0~�9�$���>�����1X��M�?�_�w�a��a�;��1%�"��dTmϭ�����w������r�b�GJ���46� �b�<�N�MnΩt��*ݧ���ܤ�bSPĵ	HB*���fiJ@��\����X��d*��d��j����˥��ݰ�ޭj�]��4�sF�u�Y�;���Q;�7��]o����f���5�X��.����ĉz�慟g��dC)��O��I99u�v�pBj넂hB�E1I�*$ms�Q���mZe��|�	��;1�s���b�Bbu�EҵnB��۩�#H��=��EL��P�3Q��wa�q*䘔�����	���7��ޔ�\}�1�DNq�j��R�yt�yH���ST��N�cN7�3knI �u�o9�.�n�Y:lN� ��K�[T�YCK�gf\���KYjR^&����q�FR��ddZn�YL�&y�$��%�[W����V�K��[��B��e����ncC�Yv��7��@�_#nTt��ܴ�gm��Z% mF���F�u�ܟ�L��,��x�u�G+��"~�ՑtL;2��ul��miԕ�[x"<(\M1"B�Ӊ�Q�r��b��~�qk�0�����QT��N�������o-S�cS���ȵjX�D����;�f3V�:��ca�=��b��3��v蠨��*�#v��Z�&����hCF�]����R�i���Z�g-G̯+x�)���~��#�=ˌ>"�鳜	
��pI�h�哫�K�<�Y>��N<z}�>/�!�!2��̇��2
j�Tk{ۇ*�h��3f��-�Z�Q]11���C߃������ק�P�q��`�l�뾠O��y+[�@�Ҭ�t��6�TF8"E�o�=�8�/�/�/K��<���g���/v�Wnn�\��5j�H����՗f]��߾A�G������]�T�3��G=����A��{V\��uh-�:��'�q�$��Z��ۚ�F�;[�u�joR�9c����R��mk8�Fu�13RM<ҍF*��7{ɠ�n}�y�DX1����2�	8��̍�)���������8`��(ݨ2[���I�+����Ri����R��� v
�����%����U] �>��X�d�8:�"�s��g�n(�K6m��;��Mn��n��Q.�ھ���>h��;��M(�z����2�l�]��ڥ���K�sb�cv�4�̫9jj�#+A:֊�7����Y�i��U��Z����������"!qWA��g����nl:	8{�*7�tۚ�-�q!�9���q����x�3C�v#��_<+�j_����F�v3�qE�(e�q�g<ob�`>@3(!�]�֌<�03ɨ�J�g��`�s'��s* ��T�`�S�����;)��	����B�=^���F˘��j"�R,8�;�u�E�k��BK޷u��Y�W7�<�<��U"3}&����8�w��<U�<~��w��uDi5���v(�H����Z�샴�s�;�����}$�A\q����e����j8��j��&������|�j`�W[����iP��3��T|xTb�G�6�c�����uP16P�X�.�b�a�uMv
N�Ul7i?��,��3����W�(㣶���ES��-LL����i�.� �.��9�V	��F�l6]�?-M�J<~���G֮�>�=��d�r�q�D�?�>�|��*��Y^�;���eCLS�Ch;<;�KT�,Ա�=6
�y��*W�*�8P^�$�O;G|�e�T� j�l���r֞�9��T�z��������[��s���R�4�h�qr;:���F��p�G8BA�U1�O?����}n������n��@?Z��!���o�Y��@�1H�32²Ӌ�׵]�=���@PG��dRf�>雉[�KGL:|dU��g9��-�zfY}����H*���7/B@�РMGv���;�ʯ�������_�����i����>�K����>�sR��]P���a��pԭԡ�1�I�뀭�>�)��<���jn���-|����x�-(�!B�ԛF��t��V`F�K��$l��yѼ��¶����Γ��ǆ�9he*&�3$��D�e̢k���m�\Ո8�6�M���^e<���.T�hd�+�8USגI$�H�rBC���n�s���Sb��⦤`�GV�'k+����(�dٴ�vɋk��tue2��n����c)+mk���Ƨ�����5��͂���E��A�S-�&�-����d�P���B\Īu�`�M�M,Ga�Jm�J�Vڍ3]�-�/�E�P=�/a�/�v~���c��\A��7*;qzq��(���0�E����t%�l�n��J�FX�Y����d�3��/�=۹�ֶ�,��B(���D�'CW�-���8��Eذ�3�g��U�t�)k�(���M�+��tDS>K�k������V���i.]@�,%`��d4�nY0k]M��*tr|(�7g['N[�4��}�j�z�Y���^�P��n��PHE�0VT��z�h]P7O�"w+�]�v/�c�̚%��#�E,l��_�[�_5��������W�An	��i@��Q�eЬ���Th�k���|��Wp�v�&����`e%��Mr�!��P����m�|����ŕ�g0(�y��u�R' ��>��,��g�_��r�~!�h��KX�~S�-��s_��y<-�9��Y�9/F�ovS��^Dng��Y{�*�Ǉ�;�u��,3�̷J���2��Ul��KX^=X&�viӊ���Q?��d	�_Qw�r�츒��p��+!�U ˎȨѤ�u�B4/����0��b��j�P?�Am��~�׵��	��)7x���i�Cz�\X]�Hܜ��)E��lN�)9M�O�D{�<����=wC�ސ̛h&� �_TBeO6�i�A�n��oS�}w
|�%A�5��SX�kԺ66]�p%�U���g�O:��l��7q��. \T$��rĕ�h�H'�r�q�s�A���Gޮ˟/W�K�zs�$�'�r%"N��~zw $ꌋ �5�RZ2�kznfg�U�u��};�>����rv'R�$�,8�>R:s~��`�3��:I����}X�?	�xI���T V,ﮒVqh��͋�YO�+,�=���G�(qp9����,a6��(h-X"xg�ga/$�j�����cl�l��T�P$	b�����},ǆ2┞���<ʊ�cD����]��]4Q������K'G1��Nr���G"�Ů{qW�"7K�R�bڿ
 �f���`�(�����4�G�*:����^����:��"���΋��֟�i�B�_�޼��'(
��7	N��@�h��A��
c��H���
�ԏI�&#=��V-[uZ�O�U�e;���=���LHh�uB	 �r|���0e4{��>w�nr#�i���u��
�6p��}ѣ�� L5|����QH)�B���@������_Cle�q�&��2��*j�����$u=��fP�xxOy|�]NE�6�	�v4o��Y�M6	���O�o��Q`-�/W�ߊ��'�!#-�m�{Mau2����#bّ��(`S������a|������JOD+�r��/��k7��z4 �5��m�i�3�j�u��{J�K�Ҭq���Ż+� ���W�]!����گ�WJR���腽xG���n�H�W�� @�1��b�#��4 ��S�h0	���8a{����U<|;�6��NK`�i�=����G��>l߇�G>�z��ªX[M<�GP?�t5aμ�f��>zA8�~z= ST�3���ڂ���q�k�i��@oF¾�c{�R�㝥�k�k(+�)wQ�ʧh��e�U_�Pe<-�j���a �̚|�Z3-c�!�gϟW���F�� VEE���V���$7����H�J�,v��d׭HA��S.� ��+�}+�E#L:�T�D�&��ꛉ�֋1���-��ǌ~�~Mve��V��h݀����h�A˰Q�m��aC@�����୵e�s�oi��hB+��ļq�y��8T3u�� �8,��S��2Ͻ�{��aE	Ǫ̛F-A��<z`�E����I�jgP#�4'��+�%=��Y)S����1�_c��{J��?��mFP: {�YK�����TӎG5�G��@f�b��w@�[ޣb�{=">ۀ1�L;.�JqI(�zؚ@��u����amd� �)�D=�)�6V{���^�=�GA����u�e��}Ea�9��ɀ��X�ˉ���P����i\&8��;皋�z�
�y5T��h���8хN�.z�׻+�
�JۺWm�H�;s�q��~�_kB�_p����V* :3JV5��/)j���h^|fd���� 3̞����<&)��K^�|�ݞ�G�B7Ӎ�}kNv5����� �lM�iG;ە�9�$(�[�P��9�4#����W���:�^���M⥂��X5��̐���{/^�`��K���܂������y���x�m�f����xx�W���P��쮐\+b�����w�muSm�k�������z�z��\�ؗ����Z��o`�ݚM|ͩ��?K��Fg.����sGg|��I#K�ey޼�NSPsw�A�(��QU���bJ\sW�@���Uν��Nt�d;��}�8��}�N�TSukn���c����|�L]�3��B�����sZS�� �Ͻ<z�)|�z���w��D�!������wVF�u�4h���R�����.m�/��{���lޚYOۏ�}�,��t�S�:1�����v;w��z%�9���+ӏ��x��v��X2�ܬq
���kC;�>En�
��m��v(��[<s����,��eyz��]�Y��	����~�����         �   :)�7/m�����ƚ&l��"�
e��"Ca�ݵ�F�Z%�P�7j�X���9�6]�"��i-b��wR�Mv#���q�Y��ډj���PH���j[5�΄k]����.1t���*L�څص%����HݠM��qZ	�6�[]-0A��ԛd�]�V�ݵ�J��٢u�r:b���)`�Yu�Еr]rת��њ0&jǨ\׬`�P,�	]����3�J�������'�L�6�;`[.��fef�[����X�\� �v�a��H���S��])�f�l�(m�m�d$tA�T�p�Fī-���%MKX����G]j�P�ZYj�7lRݴX�p�lD�V���Y[���W��ӣ�6�{Bh΍�zs��I/k�aS�(�*b��n��[�&O9��iȎI�^���^B$��]%�%6�h��u̻bكAj�-ȫ�k��af]���cX��m1a�e���-s���֮��{m�m��[6��iVNN��ƽ�T��.���HMLl��Z-"n�2Ǔ�.����m���f�%�ۖ�j��B�i.��e]\H69���1��=�[M8��
�A{��1G�E�п.���� 	pCL�ZI�/��K79���:XGdasqTZ��SD�
49�T.12&�����K�,e�-���ژ��Yt�}|���vL8:�Uyޔo:�뵳/T��o[��n�b��n �GB��0:х��.b���Gg���<T�Z��4-|v3��%|o���	�5��q+<:�¨h�/TP�5��_�V%$���c�L?(B/���������2:��s�]����3�v5o���? <'��1����>� �W�4���S���6��B�~};o����ty`:��u�4��53v�)%S�D�v}���w y���)ċl}Wz����r���
��7\o�ޣ�&)����כ�3͝�Ny�t��oz�E����UE9�!F�W�#�m�J�{��׭��?��߱�Ր�5 �Bm�}�q����1�.R���>���q"3��g��n׻�!�E`į��
�l��#�v��~�;�P#M+��������N�D�@-)cU{��Xs��v�Qڧ�uO �� �(�f{��CX��;8ۑ�Yӗ��a�릮�HZ֩HE$�4� ��U���i<2�(�O���\� ��_)�϶B	�0��(S�_)Z��mEӜ`6Ҟ�߻��~z���j�Yah�f�u�!7�\[*j�5�ȣ���I#��#y*�!jHV���%v�V ���'0�$H�w&��� DJ��TO>�g-���N���l4�cش�m-��_Q���g�qR�n�8+}��#�����T�+�}}����������M��]�����<�[h��]�|<X%$ �6	��:��P�6H���<�U>},�2Bt�`�� l*5 ��_�*�"��d��E�{�/*��)�#ǰ�A}��ҙ>�aQT����T�>��|'��*��'Z,�P�Z�!M��?/���L��	���8kBd������\�zaJ���b�cVP���p��7vy#���g���&4ƈ7��x�N�;�a�m|Aץ�_����� E�G�3@5��s|8|�����qr-04��~_y2��8�~��z���,�	�@`G��� ����2�'�Ȍ_b��nE�w��yN$���
6k`]�b�|��_��#��0}}ze��!*�<U�~g��Zx7�{��ɪifr[��r�r"��.#�u�L˶M����	�L�6��8��;(j��=$��T&H��t�� �+�'��@e߾{1��5��sL��`�hE��s�Qj�ǖ���(�ch��!w�\r��q��o�[�A����6��(BVx�|Vڼ�����D���H������Ո/ꃧ��wL���c��ߺ[�'(��`��:��%��`��������}N�5����g9��پ�����\�m�#�������f���W������S����U�Z��a5���0G!����0�8��<�D�	0��)�O�����@�,_&�v�'2�7�zDA�*�+���л�A蚷�ɴ�,� *[��ʐ7R.�w��H�wPgL&�sX���4h�	�]{���8��u���5�11����{���b��K�lO�n H�Ò�W�|]֩Y������1�@�J�˦�.2b�i!��܉Yv�Bb�!(RD�^����o����m�u�Fɢ���H�l:F���gV����^��E�5b��*�dw��x�R��4?Z߄�f�{l�u�ɽ*��ޞ�`m��?Q}<g�(��B?-XEX�ڡr�M�|��0��}y�!T�~��̬<��N�;��9�f�1�Rl�j�ڲ���a_K�ܴ������i��B��Í��<������4@g�0$�#U}4���f���cv0~ϔT��Dgdo�Kk���j=w�� �"�<|���z�J<N�P�$�D�
d�#��Xf�Y^��M��<@���ݝ={�֢yi�Z:u�a
l::�^�cg3�]Yb`tL��1���2�"Pl0A6j(��E��^��
�+ϩΝf��wq?�(�,�T�P����N֋�(d��Z6��
5��`a�Q�<`�`ڀ��ZA�[
�d�i�tN�2߾�r�΅E � �ٕ�Y��q���m���kt#�|��|l��|3��{+��X��MJ/�:j�t��B��"X��42�-�c]%n�3�&v�3i��_�
� VY8|�ȋq�h�XЮ8���{dYw9��VD	�l-��Y��//��z!�FC	c�H Z�dX>yg��U���_�y��T�[g��a���܋@���V֣�Z�!�;8-�=kHOE�ONzڻ��zV��U>��aϮr��s�(EVn^�j�A-2�&�6Ҟ�(q���n�!�ݰ�o�L�]�E}��/y_��z����傃Bo�M�>��Y�8T���>�1�qc)2NG�yޠ)f�MP<
,Lg�8�H辫pT]��&�>��FGgGO�ڥf��'�)0a���E��d@��0 G�`����bӄf�r� v��=��3�:�f	T�'�$�LK�'̿���y�ϕ[j�$
F�o��#��{��nx�e��jaăh	T�$�EKN� ���B]�j��/4���R�'��X�C*�� �޾�k�oפiڭ�2�23]=~���Չ�	��:W������>Ϸ� %��C�*���-rm�v.�l�˭��6�t�f!r)�Q46����,%�LmUt2������LBKJ�]��n�	�si`���6�]f�t@��ҷR���-ɶcl�Tű6ش��j��1��E���3h�X7]x�R��k��A*����p������?3ʋ���ȁ=�/��VoZ�d>}�i	�3�,��0I$d��D�&f���%mJaj�NK�E/qB)Ό���^�H��E��1h/JL�f�Z��i����-���F����P#�3)�s����}ޕ����A{�Uc��}y������� �^s(�_B�8�mA��P�:�m0�w�6�Z��N�_6�0�[s�ԣ-{�y%�R$R%�n������Q�`�`�mJpݵ4�u�]55�-�eH<F/F�(7t�Q	"Y�:f��K����la�=>�`�@��)����G���EF"�H�P�Z`t-�)�`B�����1���[`��R�Г�)7�O��`*C�e��3Y��@���㽭oS+����L�4�4��cr1������ь���q��%�}����0�H�+ 7�|���FYHֺ�vU+�f��n&��o�ۏ*yS΢�����:�6�~JR�cG\���N	��!�=6��Q  �=��c.)��b��u���>ּ;�ȵk0NB�c�~6��/gԊE-�y
���!��Ͽ�i�|_�o�n�,W�ޜ2���U7�"���R釻�?Q9�+>�|�M٢�r5�حm(���u�ˍ�z��h��Mۀ���+y#`zm���`(b�����s2]0�n k_F��䍠林5ɍ�e3���Qi�h O�w�w��O|�5I5�-��`�K̌�����4|,ML0�>��nH(P�C_ C�Mu����Ɲ�EHm�T�yf��ݍN�U���q���hL�+�ykܡv��ʶ<�)Q)R�I�c`��庋�t�H�^�T*J����Úan�}Q�֧1�]����I�J�Նu��
5v����$�?o{w������E`ze��s�!��u�sFs��TX5���^����0��Z䨁���ˬ5Ģ#�����X6b�4�����+B����/.:>�����m��<��O�w�U���E_�����u_zs�k1�LjF� E���NYHҌ���/s�着(�0[e���t'�|�ﵕv�?����֌T`Ј}&�P���������=�Eh�A��-47��`��
۶�`F����wX^���}��5� E.��u���Q8ՈF����l5�z���L#a>qV�1�*{.���p��?��yo��$������p��v������w��x6ǂ����@]T�V������Un�����05�Qct�u�e7O��/�u�M�椂{����`:i��u~&6��ϳ��Z�R�؅�h��V�>��9��O�G�G��T|ߪ>�\h�i�t�Zǣ����|%�&�#R=8Q�E�g��PF a�TY�L���itכɥ]�P�T\���QAw�TR�+�/� ��$�xW��p�:�>��bJ��HCC]�G���t�6�ƀ:�䆅g��n����3L3�� �375m�(M�B��������a�DQƆ�m�˜�s�;����ơ��]�qik��m1y���E��@��gL�����D�D3��aD^o�|0nE���Mg:����W�q�Ԝx�G�G�C�li�>�v|���xe�9j�qC#�m�1�a��T����7�>o���ñ&��wm2�,�E;呴_�3b�z[$}����!X � ��,N_I��^� ��=Qa\ ��JBGUS%�'s9flGm�UG�/��r
�AX�ת�m�&�*@ @!��H�ݺu"��>h��0w���,@ϰ���x}v"'"�H�'RaQ<i��� ���$@��[%��Jj�E$�;����߈Ͷj��<'���A��E���ι�;_��a���aG֘_rh�Ǚ��l��
aJ�m�k>ƠK;��,�I9���0'�L����Y�|�GocAm�ߧ]:WUHRE�䇊Q����&`F��P��(i�|.��=><R0lv27�&�7�F�z�����H�\��{A���c�q�ز�Pڍȫ���D����2�����Na΍��� bx\v��U�}��P8[|#��!�[��yg)5����L@[|�g� ���  =*' z���;�R�M�D>�8u�`SVW��j�g����B�#J�������h�<�b�ȅ��h�Lњ�޸����(�x�9���Ey]�4����� ><K{��ci ��*��v��Q ���U�|��`�£P�t�ua�$�M��j�DA��x�jWn--�4�8&�d�%)30�Wu���J8���)�<�4̽gC� y��Ր#��ˎ��mv�\�
�r�dQQi`��� �!n����ɨ۵���5=���V���Q@�����0~����b"�T �y:� �5v�>�,��]��M~(b��lω�C�b|i��	��}*�2�Q�8���+F�O��BO����{����L���N;ݏ���GZ�$h_n�}�;�$}�}>@ �I9�e��,+�6a���-ҺГX%����6r�m�{]��t��Dz4�6�V5��ư��5�kUe6��Ֆ�.�	�]����˗;s�-7�mN+^�sLd��m.�uJ�{9����2�Ԑ�c]��l��u�n��c��Vݦt�����
>3�AE
�}y��S���
iVȬV��������܀U�gK��V})n�
><Y!b`��ry69RVr����r�ʘDY__�{����j�H���L�G��X���`���D!=���I���)?0t�;Ÿ����
��g(�(U��i;��uk�ka�՗�a����э��t��%��8"?}�Qr���A޸��ޭ{ዤ�u����T�h�3�����j����q�~��\(/�(���H����E]�a�$�$]��|Dn�֟ 0N�>آ�*mTȣm�31�Ͼ�'� T��[�G�G;:���=�OZ!g�B(~"��ўF\-��h(�����m,j�u��H*,��Z�|[�ρ��ޓ��J�ɒ|\|ы� X+=�J(����)�$�P�Q�$Үl񪫛U�ԏQ���ݵ��v�=�nXֳOn�W]Xj��>�ݲ��@�g����w�."������IO�Y���&�M�l��(���l���]
��!4G����_[�.�W�ϭVb��x��b�	�� H��QZQ%+�od3\��!��JTc��Ɓ�[��5��%p��R���^+�p\)���d)f�^�͹�mc�k�w���� �3;l��FR *lC6�/�ّ`�s�X�h(`�y]w��g��]߳��{����@
�i�d��2:(��g�{.����fV�KSL	L|��}��G�8=]LܠV'��#mh�k�$�M������u&bY�w�M`�#������L�v������b�:�
6w�� 	�������%'��(` �.�|���u��!Yw�ޮ�zT�Ό��si�8�����*6�!j�B�mtc��m�Dm��;i�~���f.��W4Fb��91�}.P,כ掇�+	B |bQg7���>��� @>}��������XxXDō�7Kh���1V4Na��\Yj���|!�C�P<|�6�%5BjlUN��d�*=_}��)��Z`��w���Ϗ��*�0���Υ�y�j��,��8��<����mS5@��?x�T�U�y�g��X�g$Z��Z��,bѯk�I��Ɏ&{rQ�7�-։���}~I�-,H�����Q��a$z�kE��.��#��?R@Q���Y' 'm3���)�FQ�a�%��Sh81��x�Ų}%�]���*�0�Y`�=�m�kF�q�L����*j�롧Y�=�I��B|�U=�����E��j��{�"�����轾���,}~VX����{��q~pU��/�Z���c�oi�:+H]��2828?wY_vג�tY�8^`���B������B�ܾN����{��^�=��CT�B��Ls3o.�ε��J�8R�v��U,ӻ��k#'mv`�������F��#�>���l������
Y2��^�c5�mmx8�c����9tK��NN�U��$�5�����3�]޹zZ�l�9��'޴N���-<�<�+G+��5wr.v�}{}�os9���E�jR�E������L�'+�Eš5���y+����������XŪ�ɱ�[}w�$�Wu��?�g7��H��ю�V{�	ZDU��v�?>A�|.���|��C|ؠ~\�i/~/��2�O[D~c�7��]��GCG+�ѹ�� 8c�y睹�*�>�,���ʊ���>n<,��j���b���֜A�E.�>ǅ�M9���V������GN�L'��~����@��Э�W�s��Ha��[�f���.��e�A!�RW��}���ڽ)C��H,���YO~c��
i�N3\��c;4���4�ɦ1�#�)����:����A!T�Ԛiu�[D���8f��E�ڮw�z�:^��.R\��9e���s��X�N�D���1:1�QD���J��s��6D6Y֠����Z�1��,g��|��O$�A�b��]ƺ��)6�f��߾k^�W��
9���j�\z�PbT'v�+�"f[R0�5ȏK�ج�q
S�Gv��L��.խ��L�� -����] h�M��yV����F�9h���}�Z&��	ͯ����\�G��`���;�uuK����*��
��V<�D�8M�D��E r��eJw�hmx�Kǋ	 V3�E��8��h4�������yKt����"��O6rT5շs��7�����ӄ�J�<; ���6; ���'G��`�{^%F�����vP W��l�=2G
��b (/�ݴ�w��#�m���|�A��nRۘ=1�|E$N�:C�2�H!�\z��Ϻ�Gse��c�eS ��h�^����9��
�P��h�Yfu���l�h[��ch����4oG�X�j�R� � ���t#���a;��X���r�Qۉ��C�;�B�7F���F ���U��I����(��b@����=Ox�&�bA|�!�t��(�qkoH(+,�������P�6]���/�B�Nu�| �<��*Y؂u*����]���ݨgoB5}f�4�$G������$�ݘA)�{#�H}�A��=/��0d*:�Y0��O����U�wmK�>!WST}�=~�� ��TI�L�L��U}�Pѣ���$]�@��T?�%;zE@6�[k�ͧ���r�	�cey������[���h%���0�|ǳ��٧݁��Lt��g���F���������^ґ�	}�.��b�6� ���dJ��#ՖϚ}��ǚ�!=6�]��S��b*<����K��E^�<��;f�6�}v�|�<�WJs�;�9x[�4�����p K�^�WI5��N�J��FŖ�����ڳ
Z �(�����*����k��+5���\/,�y2K	$���.�-�H�1ŷs1h�0iX���,SdT؁Y(�ۈ�.��mY�iv�������]bs���Sk])������LKH�#@��?	Dh�����L�~f;���lO_(Q6@+��0�f=�����׻�U+B`Bf�Z2�p�J�����L\E�t�����Hڂy�^�(�IeJBcxj�~�<����Q�����9PCeÞ��'�^5h��_�:x���'M��ܰ4Xu�<�EwhPp)ݍ��IP��=��������9���Ң[k�p"(�h�#���&
��1����4�`����,��(r���9��}�ǷW�ҀVq�4��R!�/!aK�T�V�\ve1̫��hB��Ta��!�qiuL2�&3��f�ڡ�جn�}�@��Y�����qe4���)}�}gew�P��`�m*L��4�*�s13��+ز���W�U�h��M]����B>��Sc����Ω��Ӊ�S�൰�������&t�W�a7��7�	���puIƢ��b��[nj�m!fE�k��b���iϯ�Y�q:i�F"���#�8��P��)��ﲊw]_z��k���q�ʀ���tYB���� �]ͨ�P2Z���O!���ly���-\��}5U^s��4�D3i���yL寬�]YP��+���tcL�'��]��Q�8Us>=�鴾�auh���:H^�-���j�{�sS���D�q�S���[�붲��!�cP���RJB����Qd��oK�z�0䉬<X�W{�g���s���+U�6[^���5b!e�� �z�ͬ�v�<*3�9�_e �-1f=��:E�}l��!��/��|h��8�87�����U՜:�s���|]s��g���χw� ������wԾ����6b��}mKl��`���|�[��!�	岉���u�lz_���{Y=�ϝ�4�ԟT�Xp��>4h��yq�i���\	h�i�I^k��%��( I�}h%(�x���+���f�v���Y�i�z�l�AG��U�zh����hg�����"�^ȫ�+ mG⬳��o.���8�U���ob�r�"�$�B�9B��A�4�b�"�� f�GH�j����f�0k���_O�s�mUҏ��{�w"������ʘa������#w�젯�Q$�N���q �&��˧bm��j������p�馘�����|�I����ێ�$>�����uziĝ�����\']���߰V&���gWMT^[��u�x0p�6�|廑��A�ՆyJ��Qf��-�=�q���n����<�\9�/�ø[�q�K?���1�J <�=W��~(#��q��[|E�`�H�c�m��^��3pu�e�Ύ��x�� �d
�|������(�Q�%
~q�LU��8�5 ���N�{�K6x�i\P�L�~i�/�YvI��l��p��p� �r�@� e��:���ߒ�
04�Ԥ�բ�Қ�[�Ζ��)�۬-�i��O�}�XY�9}��W5τ�����m}ߔ�9��[G\!���ػ�_G�#�r�J��F�,��9���^Eb���nT�O�'��������w��>�E
;�`�_6���Ys��W��ܐj<+��ъ[���o�tzV�o�k�}q`�lh1��d�O��2���Η�;xT.�«��=N5���!�m��hWnc^���:ޗ��A���S5�Kݗ�0��S�<_^^�>mFLW�����`���� (F5�B��9�h�DqŊm���4G��g�V���[��E��u�_����뢆uT`��㸢
O��f�2�ԗ�}�y2&����&%��6�>�{�k:��o.d����b�|>r��:�oPFu� ds�G��/Z� �X���0k_E�$�&�]�ie;B�A����%�g'�yk��>���F�A�2�*8��qַ��ȫ�*:N�s�ը��OR ��s�뤁\i&�ƍ��0��6f�m5�l:͘]�e��َ �z>	B@[�v�>i���jݤ��\a�_27�cf4H�������%��v)����6����B�����Q�m	�KXt]����Em� � -jN�����H�L��b��K�R��:1�"�uUF�w����>+�ӟvLL]}��W�%�D������Zb���S`�U:�5K�r���Goz;Hx�D�-m�ٹF�a�'*>+���K�� ZA�^^l�4ek�;T��q��<�oCN5c����an��@��� �eO���[Zr�#�knȧ��{m���H�G����d��%տ�(�k�O=�m$��xq*��R�+�k:�_v ���U�X��0(k.�Z��C	 ���۩�a�K�c���5��vw:�L�\w'Ez2���i���װ�q�}�*��I$��$2M��ka�:��f�u =�a��j�x�1�U�*��j��3l,\U���1�ed5V�I�Ѳ��.�Pͱ*ѭ�gfkz��8��ޓ�]5j��pci���-�W�i�Vx��*lk�=y���ye��v�<�M!f�R;\�ջE��H�/�2�7���W�Q	���NH�����tnRk
'-CϖuN���D���E��`UZ��-[�zwr���J���a���6��C�u����,u�a.=�L0�&Y�7IH��TF�*�6�;�;���5B���a�+��馶�ܻ��&~�Zv�a���Qn&j��we��:�Ո-|�,:�ա|����K0�c���W{���I�?�s)HԄ���`N4QeT)��Ue���I�C���E
��ä,��Z�>򫎜)��OqR�ܳ ���I�����J�[p�m��䝩����P;6R�2�h�`�W��}�Β����c�T/�������B8�X������2�(n/���#7�=*�"���b�����/.��q�������@�����W�pv);�={�~�>�r��]�9`�V�M|�V�q�7�H�>�	^�&��M�@/R3MIQ4ń;%�h��r��27�n�g[.-��AO�����t}^rx��9���2�TL��m.����ݣx��@�tC���_�lO���=&(�l1�uWX��|v�F��V�dp�����Q��T�	!hG��#+ Oz�.S(R�m���u1SDW�!�vfwn('��6-`�k6���ę���A����K�I�D�'g�B�ؼߩ�Ʈ�d%��3�L���Դ2�'\�A�`̧c:�I"p2�8���<d��ث���,z󦬓>Q�ti��O�غ�)��Y�Ρ�m��@�eev�@ 3RڔLڼ)ݔ@W�4��	l)���X�oxuN�)��g>��4��.�4��2��V���_���87��9[�!+�p�ͳ�K%kPb����HF���Hj�w���T��f :���@��sG�\b�,�p��N@2���_QF����zB���Y}��ά�v� �e�Ga?��UO�LV��>W�/]*�����횚V�ŭ,q�qu��d�W]qy+�K���侙{�!B.��Ҍ5K�Dw?��i��ޱQ�}b�x��U	��$l���d)%G)�,�,��z��kɺ�fNtj>9I�D�����xhօѲw��`�R�|YѐD%ad��Zg3%�OBX#dJB�^��Ds�e�2������Mg�b�qs��th��)�0v�]|NG]�3�@����g1�[}�1��E�\C&k�*��U�w+8,\L{��ZPt5��+�i���<)�616�C�U[TǛ�#�u~�Kai�	�
��ת��yt9+TG+;��|�p�0r
�]˹/߃�}�pݲ��K*���L�1�a�nX�i�͓]Ϟ���J	=o�"z8~Ѱt��@���Ͷ.b]ֺ�i�� ��`��+P���m�d�-@c/4���٘T�B��A*�e&���dt�6�E*�e�5W���x���B0�n�!��d�� �3�E��(��l��J�b2]ʽ�1a?NR<�ȾB=���!���Y�eb~���ǂ�F�OzTaR��\�����.z�b�+�"To�2��T0G���Gt�o���t5���Z=�b��ʥ�bjɗ�X+ Q���rs���M�?��پ�u���!/3]�[;ϯCȆ�����~�UG�ճ<ìe��k�|���r�sbcc�c�d\FA-�U	�x/�}������������BW��.x��ݤ�����
�ƫ>]����l�����O۬��SS8�r��&{	Ȼj�+�o/ӌPG�c|�ݗ<zm�:W���w�W��\溼��.�I�Yg��j��b�;��<������=��ކxi�ڭ�ݬ���}&�U��i��ɘ��I�r��!��!���7-�\[�N�}Οw>_j��J}�V�;a;���v�G��Zu�_��1��}�eX�ұO3@Qz��$�7v��������Yڮ��짳{n;?=�㛜�I�]G�|�����'��O	���{r)8n��S��������u$�I$�I$�       �   2w[cuI�j)������΃���cE�4����Yh���Of�6�f�f�z�1[��TĨQ�0������R�n��pK/H��vZ���Q�[ն�S76)Q���n�m�ׯi*h�%�Y�Z6=c\�����nj�u�.��I���l���ڔ�l��p��[�W)1b��e�h6����i����ݭ���YfE�4u�!j��GR����m���z]kV��H�傺2h�Yq׭��rK�:Tn� m,����1lƁld�ܝ}��v����&^��H��'�-��i��ܭ2$�K�\L�J�(B�[A,�u���A�ٍF`�	v�0�٪kev��n��T�ڑ1H�#0�R!�i`J�+����@f6��k.`��uuIvR�44q�kJD�5����B8՘�+��Q�FvZ\�7a3u�a5ae6�����+b��$-]�\́�6.�Z\D�ۍh�[l��ar�]��*����۱m��lH�O3e�ۯ=��#c	���d^5ڛ l:T��ì����6�u�c���& �u��.�Ӧ�ݸ�1�ƃ�iA�h�͔�
�o� �G�>�/��ܒI$�B���r:���Ӝi��ʽ�{��%�nc4���u�/]�i��# �n,��[6�@��CL�,�P���a�%�K^5��Ã��s�`MJ�ce��i6٨�s`I �ےBQ$M}�{ݤ5`ꠕ�;A�+]�2m�3Z��$�"�
��߶�	�T���eayFg�wi��Y����Z�̴^�` �Xǃ:p-�3�e����U����	���	�-vR5a�X��Y1�Gl>���YB�p%i4,;eN{�7iي�.%��f-�T�4�d�!q:(�fz�\�ʵv��q��u\}���MF�Hԁ4���8l�|t6��h��n��rn>IAD� �i�0塄Uˋ��2ju��C������&�n K�٥ݕ/��mX���������?'��M{��ˊ]��	]�2u8Pz�N4JJv�ʥ�DZ���G2�TʍB�R�/a5�����"�j�rh�)m��h���7��M�+��{��u�{ ����(6�
���%���R{�H��֮���0ǽ/�J5�:��.��kko��Z_���sz�^W�,,}
�`����5(�l-a?����*vH�n�g�gC|�
��=���T
�_�����YWA�lM�O�0]�F�7�c�taq�!iq�I�6��	UcX�yϞ<�"� ;O������/�&г����2�i�
�
H(���D�G�]� ����>��oQ^�>�E*O��.iah����������[��TD%�����Iϲ4�:V�4c��6\A�܆�Cѓ]u/K���auӽb�B
_UP��\]�#����k���d�>�srh�g%;��I����� M��8��6�12N��v�pX<����K�"�bT#�1�R,�tQuH@���[�yu�3W�����%�@��.���y�7f�+���%O���C���T����PK�%���$D	�i?���7�˯WK��ӣ��ٻVmq�kF(Yc�A`�F�Us'��^me�8��+7&!J&�s��� ���}
���7�S<�1��D#�䭽/�k�H&Zj�� �XKL�&�&DtrËŃ���-��LU��C�gG��}�w��{��Ii���{������|�ht܍ڹv�8�Tz@�R<צXf&H����.�����آzn�\-�-��o�"bRY�
���zp�#'�v���ҧ�J�����4��B��ED����tpN=\c�w��(��w��BY�9F
��Ԡ�{�}���=�=9�v�

R��Wh�3�Srp}Yܦ���$���y��M&$l�fɗ/ޢ[J����f+l7�]�_� |
K��(Q;�{�vS��$��	+�xl��t�AJ�֡jjF��Sj@��WYV0�n��ΩM���k��4�c<NI��7n�jX�ą=�&���Tf4I."�yOH���^�x�y���}ȿI�Gu��ȷx���7d����?M�H%N��J�ϹJ�H܌�b�4osh*k�4@�l����L������|�������V�G7�؝eS����#5�L�D����;jvHx��)��G�@�<�j+�m�cY�i���r"����(P��Ni�j�0IP@B�)�P�*�b�"����2�B���S�7��ʄ ��+��#6�S�����a�c�%��"\wb�9���N�VV�����h�K�W�I$�H��JM��b-�^+�!fa���ͣ�&��o0m�b�&r�%�nc�*�1lc����(��]��"�%v.��XJKYej��Kk�D�)��Y�8,�\�G8�Vb�z��I�e�Cq}�)ξκ�/6u�XP� a�P5NHm�
�feCZ�Q�|;a^��BF���]����� }�s�))�j�S�@c�6�RD�[nmG���(<:ť2�6k�%�5Ic�ʝ�Ś0 �b*w�Tc��Ão�`����E� �É����������Dq��s}`�S��;���������%��^^�zD2�3��J�!�{
ZQcf<Ӆ��OVQd��2!g�	Ɠ�L���M��̸#6���v�`������b�I�2D����[�U4;|��/۬���%����j��7I$��W�NV�휋�\_t����{>i����E���ҎVM��@fw3M�G�t��j�)\#�.����ˏ���}��7�ߩ��R����FT�kG7��E|eɾ�1���(jS0�3[�ٽ�����lz�/b��"aDW���A_%�'�~�u����RΓ_�VBM,�2�u�ȧt�t�4�K�)��x��.+��ޅǍ��Wj(���gm��ո�X�Ɩ��+��9�*�2���A�+2&[}�3�o��?n���6=g��1���O�}7�4�6X=�t�v���Y��kHX8v��WGmm)boWNEaLR[˘��ٷ�lh�,�$t���0���$R��7��%3�H70Q��^M�@0��P;Z�E3|��:��ݧD8/�����_�=�U�):6�Y��h
D����W.�p,���l��7=�&�{sD�3��峞"�}xǝ�v�ݟB�!��߇{��j�2��]�s�����Ո��m(��s�1k��c(Ӵ���Mo���cN2u�9q]���qLK8#��bFA�`�2b���B&q�
�s�u�N���v:Ī`�UP�8���\ޓQ�6t,�ZL$�r��,jd��MU������;׽���q_WUx�ݤT�i��b�Ĕt�f������)�L�CwWS �؊ �y�0� ����X��ɯ�BD�%�^��>:� �y�v��	զ��=��,[��S�0�U�ä潨��S�lR���$�D��w
�u'�<��P�����z����/��6WT6�R�:����q�z7�ӄA���Qw�en�έ�-�yN,�>�y�N{��y�کV��A���S�MXe��҇^8�{��[��W�!�<_$8��d�{#�i٩\��6Րuj��l"�t���+`�5jem���E"
���6\ޡ��c[�A8�JisM,��}Ќ"I�+I���hP*XB'$B�:����\������s��HŲ@Hm'X�8���k�8V���7F܌5]3v��nª�0�l�Q��)EV:��i�&Pu�i �N0\d"X
���cV��r={ݨ��N45P���A�##��B���]��✃8�MI	󨘾�����r�w��z�k=�/���GN��Ւ��pŉ����Pe|!�6�"=곹E:�&7�2޴�3>5|K~�W��}p .a]'E۱,�V��Rb٥*��l�[sx�%�fL��YR��/]c��+&hJV+6�qK�-���:sZdJ��/[M6��shb��/JY�]h�[4.ؔY]��K˱�e�ѕ
��A=���J�9ƖT#4{]�p����Ռ�S[����b����S�뚣.菖P���m/_��	���\��UjXDKWK3'L�Q�Dą]7R�	�IL�Ӻ��Ť�:�@C���44� ��� }ׯw�1�l���%7)���� 6ߺQ����7�3�5�F�p��]���[iZ[�*����b��F�Fk��r߽�=���7��T����d��������hWۙ��*�8�L��3��T���noo�5&7��R�qN�\�4�L�/�X�N����,�nR X��lZѸÉe2�p([�@�b���}YU����`�l�ʻ��$H��]qܑu[��T�^����e�m6K��^f���.�T�c���ޕ�����B@)$xe漭��i7B��<��7�fs�
QL�l�̀����MPs4�\�%ҙ|�2rA������׷.�ͅ�;���s��3`��N���`�t�9 �I'j�u��{��_h�Ά�������Q���`�J��8�>��~Y�t��Z�Ike�ut�g3��'#$�\��J-�6�cŰ�t�j#.g S@0���F�&s0��6E	m�Ѳ��Rhr9T	�y���^{WuQM)�Hц<�aQ�^����'��І���b��#XРZN�7�ݪU�*n�K�tu����g,�ɢ��/��W9�<WXk%�R%��0���QC��be&VnA���~�~/��W�O>�����~���ܬ5�X�oUW_0�jꏚ�=M,1i���;�{�gN�[�@��kh���#���6��5�X�{��A�Z�c��~��R��ĸ^���f��ul~у�;�	}�^��5K��Ά�d�Y�E�s�L�E�Qbqq��m���3N��k��<�/�ž�5Ӕ��y��DNnc��ݩ"|[�V:d9�if���F�ۻu�3���1���G��E}}���t�v��y�X����ނ
��%	F,��x��	�x���T�4JA�C��g��e�3��@�A*����%&ܓ��x�(c��̿^��=<SwU�Fq��{y4��%�+`��V��')m��	�A"]Jr��Bk�Լ,�ߪ���������d�ʿ���?/���gb�ɐĢ���n�c�Z�D���Z���`��Ĥ���u.�- �3��2/i��8f�ww}9�ue�o�Y_��� H�����dcK4<�8���_vq�T���@�v��w{#ս��O���D�j#y �)N<6�&K��`E��J�
6���٪��P�p=�9{"�M�Yb�̍��6��v*ߒ �JE{�`m�Dؒ��[b˅WI�˽�l�P�a�<^�v��^����QG���"�p���v�e]=���8�K<!P��ٕ�/���������tBv��J�P7I!QJ!險��9����j���uض�
��z8�l۞Z�|Q����	�;A���h���l�+`;הէ����~�e	���h&҅M���yuX��K��o�-Lwv��Y�D����[f�1^P�-�cv�"�e��h���D]y.���[�&��Yak��ت}��Z\t�1 3��Υ]x֋q;1����KCxk��Hi�q��7�a�4bSh�UӰ^X��dz��S�3Ok����Б@�I+�b��w~���kU��'>h!��t��O��H����R�ݨ�U�ld7�K���UU*1w%�C��c9����Q���,I%�xX]2�.�@���z�|ZG�Rp�&sS]�>�@x�m�a��K��$s	J�3lf���:[��f��&si=
��X�m�Sα��sgY�ܒI$�D�=�k��Y��b�0��Xn`�5�oY�7Cu��j'L��\�]��յF�p��Dr[��W`�X��f�ԗLF��G��5�.�Ivf��͊��b	c�ѷP�łJm�#�ġ+�۪�H��9]�^u�v�#������ "Cd'ș�ۻ��;6���;c��KO�_n��	����8�K�|S
@�7QE�}�\��G����4�U��}��;"W��l[���޽�A�{��oQIvkj��N�Y�������c��H\hq���j.�i��%!�Ùu�����}�͆��A�&��;|��{���7hȻ�yk�逤�������!:�tۨy5aԘ��l��V�+�G�������y�.�؛M���,�k�.p)�j�t��'�1�=�:���$�:���gD��Th�)��FL��s�A�W�0��;�j��6#����K�f���a�ن����lf�W�!�m<73���	�$�\7�s�Z�{2�j��u?���@�<�	����J����ʅ����u���Wp.#b��vg^�V�D�&C��W��-J���7:�1u�VqQ����'�X��ƭ�Ues8��^1	��t����a�(M������o�wؑ�pq{5�5�r��d���v)�vW%����M�AA#�\���lƩy����f�በ��mu�Y�.���l�4���]�!�Aֆ���{.:z�DD�ȕ��e����
�]-�5O̻�͙��^��ǆ-�C9��|��+K�DuUK���T��n�PWw�1�!��R�AxIۤ��/��ð{�9�_Y�P����f��]ev>����+����C����h#�D��TTC���RoA(�#��=�'L�l�}��ǉ/��'�ט$^+V���c=w��S>���0����a�{��6|�a#j��A�*�6-۶]�Y������U�Gx]�2BB�4$�Y�[��(�Ė�`���!Z~�f��ޞ��E��>��49|��J�dM��e���(s��L�q��Uy�D|_U��U@����
 ��ͷ��N;B	�̓I��L�b��İ�t�E�I�g{��y��2Hyt�(�[�r,(ؼ�����px�N��q��AH�9����k�0i��m�a���&��?&���٭5��צ�mWS�1枙���v��[��}C�eJe֊�T�Λb���R��*�G�q�`��e�vvlAL4u���5��z�^S�,���B���s^N�v:,(��8S��j���^�ݔ���ؼ.�D�j<$6�x�;��RO6��[�4�4�5{�-�tr{gP�G��djiFb�Z�M�)%W�TQD�1����RȰѾz\iU�7����],؁�c7��^dRmy^.�a�ZV(n���
9�SR��I:+B��mr�]��"-&o��E.�ٱ�dh��M�z�o�Z��X���1e�Ay��>;�Xb��M6�4RtE�s(C2�S
P�ym+i#��pN�UP8��L�d��wS�E��eB\�>�]���پ��=�$\�D�����֙� \��}�e�3xuS8���jF���nl�H`в�i��닜:3V�\�g^�;@�P��糳�#n�79ƴ3M4 z˘�m�Y�n�1�����M�P^%䭚�ޖi�Wok4��\ζ[.��s�Y��jF������Z�B�M�Lh�I�W̧~]!J��h��h��KF磗�=:��/27��CN��.���G:A�!�2V��^*f"tZ�aԅ�縌U������^#\���{��P���)ޝ���Y��F�Wp�Wh7@�;w��'T��o���>_`Wi�����@�G�`���M��tR���;��g��OIE�1�{΄]uF�y�P�.��6�=-U���f����_�F��8��[ݔv��VUڤ�k���;X(�k��:�����ޡ�R����5�z!���7�	�zd�����8�֚��kF�SYU|i�rwm�<���N�F�m^Ν���^�a�ݡ��'s^!���]U��b����)�R�����)!�{�L�^�{-����ǵ�b�.����:Y{sd}�<�Nk|�|�>mڎ��k��i��p1뛇�r�����^�y�M뻰��	�Fxo�L4Aܸl�=�[*]a�w��S�(��ҝ���N'�>���m�s`ZMȜ�}w��R0ֶ�Ye�MST�&.�T�zZ�k�|�9�O�[F�90u(��.����:��.������(դ��_�1����4��HuK�:Z��o����őK�+�\^��tJ���N�u��ua#*����#�4�U�h���/��7�B�{�x���x�ڍ}�j@O/ow����d�y6�'q� �q�L�g�L�'�tKT%�0�B�C�1���;�Ǳ��i���	��Q�:�r&�E���7�T)�mm�/�LtX:"Ͳw#��|^�x.�61��M�/��lșd��10U�v
V2�W:��2")�F�����vH���V�0�$�z�9(����e��=���Hm�%����>�UN���(��i���*ɷ�_�7,5����"�AC�C?B_t��aWخ����+`޶5\=B��'M	BU	%�����r�)|2ٚ�����Y'�zn�r�j�����wcwg-���%Tn:�p��	*��!Ey݇/	��*�VG��iԺ����Iϔ����3O�Gxx��^�9�C�M�U�=8�]`�[����i��A��H�`)�ql��kz.nv��߫ZF�ܨ�P�V�p�X�ѷǖ6v���#f���K#�I��f�W��8]�I�T4ϑ!|����.�A��+d6ɴ^��Ò��dk��C�C.�e]�s=����Fh���A�b�1��1�hŕ���BRD���D;��j����w1ڷ{wu����"!ްBR&��(Q|�>;�e�g�M��������hUk�K�g��s�H	�uŌ����n�+���Tؼj��U�q�U@���h����޵ӥvP�� ���ZkoUs��Vr{R����R���w7P�|hg����dm���𽪬���%.�;)��W�N�*��0��l�My"ӊ�lg�&[��{���v��&�z�
^:����]�, _v�*[_���Q�"d���p��!�ТYF��	or`{ݢ�Z�)9$-��s�\���n�Ҿ.�;�N7ü��~��n�-�cM��F��#��J}���C���Vn��{{g�Y;J?n�y��+ ֮V���bP0Vq�~����N�W�b���<n�y�OK
��`�j�o>˥����n�k�B�kXރ;e���x��{��[�zu�;����3��q�a�Y��ͽ�
�</�I����Yڽ�+lݵ�����』�>@         .`   zcOnY�9�D��'C9a��E��x�q�k��YKJ9[���es���%����uպEfK(��y�`k2mC���)���	t{�6��R���j5�K5��O������@xIU����i�%�3 \�YH�m-�L�n=��u�u^��ł��
\%my5�Hm�v�hA6X��{v�M٦�z��Y��]4viKe�#Z4�i`�����p�ӌ��3�͔]n�]t�p6�b��G�#hԙ0�9��.��u����i�0b�gj�[nH�&�2Ո!a��֣����h�.���J��;�cfc��,�Y]�f�"�k�ͣ�z�yI[�B���L��E��\m�R1onD�mE�*���˦b�"ݬ`3�Z�!��ʉ,3��).��l*���v���mbzd�i��n�%�J�J۫��4�L�%�[X���n�eu�R�DHKZ�0�MaΎ��4�BU0rju����Uv.v��WM�1�s6If�-�����܆��D���+�KN�k�׆���6P�7N���"�)	��r�un�j81���i�`u�M	fJ���"d��e��m �E�չ�$�.�t��#t'Yz�4+�B+L�f�;F�].;6 mK�+��P�����V+t7\���C[�����U)y�����Q�`D�v�%�Ѽ-3��[]hCKF��B줳\e^Ѹ�o1Ҿ-��,6%-6�e� ���Jl)A$ل�`�iVfz�u���3󰧡��Ev�٪���O�-���"�Qi�0[���t��t#x���Gj/O	��&�!�h�t�H�&1C>w�SX��J/�S]��*Ѫē
?u�1�,����h&�Ѷ�\U�ܻ:��uQn���ٍ'"\=�h��ȥ��7
Da"A�h�#7^v%}�$^'.'��s^3%9уO���;|�5�*�[]�-�i��ˡGL��۵4�k��1���QB�1Y�!j�����ʱ3�t����O�Q�JYo>z�(o0����E���GfGy�z!�v���y�Yy�<�2?r�=��`��{�;qctlUb�
}����z6�Q%"�+���S�{���P�(^������XN��]���DXJ���]��,ְ�����Y�1
���f'_nu�k�AFT�T4 �������u|�M�;��1�r4��_>���oL�qS5̶)��.G0Ȥ�ٕ%��Z2�v�kKf��v���kj��mZO㻪,(�dG¨\nG�l0��ij���iG�E��@�l��;�gIul��(���q���۔��Am���;w��1�c=Dk�m���N<�n�k�'��VO^��_M��,��g��W�v;3u�Y�7ꡩ*Jn�6������(�٪uD����혶y�8<Ӈ�6~�GNu�ۂ-3��c��vZ]����E���� 1�,]l���W���W��Q2�E��%�����l��l�Slt��$����5e/�&>�ιw�\'x��UYs�}l>I�5��l�b��!XN{$�x�M�v��|��#4U��ӳᨬ$�����������Q��ڬG�N$��״��2�1����H�G���;�`�qVwm@l�t8R�iT\{��n�2�{s�r覇WƓi�E��[՛U\��+P#��+�"в,K�%xzI�����8/,��L��r�8�����wo���P��Sm-��Gn��%�q��]V���t)��qx���I�xpa�x6e�m�i��݅�Brl�@�Ѭb����9��Cy᛽1�f#�བ1x�EG�'���+�LY.�4�`!���/0��k#7�*wr�_
�%����n�7���p�f�j��$u�F,~:Q��������g��D���V��ѥ��	!$� kky�ö��ުg���7!�u�@���G�S�g��:���j����}/&��g��f��<�������$�Ip���f�Mo+��	9&�r¡li*�D�[��BYc��C<B�-�1Fg���n�t�s6ɫn�Te��J�]�[�6�pɸ�Y�\���ƴ�f���j,��v�h�WSM��:ǲP��v��KfԖ�@�� �&L^��C(8�P�qauU$�ǖ�i؉gS��=FS�1�`��i�3F�U�f��Xi����+.�.z�ĺ�;��m���g2_m��N}�ʔm�6atW:�P)���b��ȷ���Su��Gekn��$��6ƽeK�!�ܬL��]QR@��q^�����(�5�#�f9׺*�p���$t^-��[��RI�f�gYgk��p�됻ױJ����߾C�;bM�%*T(Y�8�M4Ҭ���k\��g�,�}�O��@�mf�T�o���\��Ъ��;�d	���J5Z���CQ��j	�����޽9���#�i=��H�����4sA��ϻf���n�F�̶��i�N�$$}v���ar�C�K�ηb���9�HCyN˱�)W:,@�g�Ϲ=��cl(�E��{Z:�r4Z����x��Wi:�]R��Rtۯ�a�Sݎ�!��a��t?����C�����4��z,���Zd{q�A����O�ixxNf��� ^���y�j6[�P\[v�nn6���ٕ�j��[���|�j�&H{���5�R��RtZsQֵ����.�}���T�@���ll��v�b�[Yp�7����7T'X:�֘���E�)jG^������|���ف:�5��ݯC+G�ñ�sm�;50�{A�y�壭��?�u-�u�T]upj�*�X�%��&�;*X"N�U�~�C�i-~�H��U%�w���Rc`t�jHA�K�p~t����1Ť%����:�[ߒ�}%k�����W�o1�(�!M����.��Y�ہJ�5]�c���`��V]z`�e����9e�G��A8��K<��%#��66����wI�����z�\�n����C�jq��tn㦤t�
�k�$2!�1�,K��U�̝x.�۶�rj�-�_Vh{���-��ǡ��h�#r_>�w����6m`�M�s_m�E�v�&�9"��9=���N5J�GD~-l:��ٚ�N �͐��*)��-!1�q�)ö��\�Uú�ݹb�f���|l���VAD� P:V��`�l̸�0L����.؛M��z���=|������R�d*����!/���r×C[ׁ����5��}��(��3r@ع�Q������� �����J4���8¡m%X́ڹ���P�� �d���'�	⻕<�3x�-�8�v�6�.Cvܪ�f�=���p���42�Ũ�7�޼=�M�
�b�
G���Q4,R1P]_,��3�N�S!�\�����rA�'گ�܏���ݪ�۹���CM[�W���ɦ�\����;RI$�KQյ�cD���
ҥ�h4\�������.����iu���L�D���siu�W5��>]o����P K.t��8��m
�.Է�]��%�2.�ĵe�2�3��ث�vm�&7 �Cl���m7\ݶ[�M.g��֥Bd)���!K��t�?n[�Y��{�ê22zY��o��QC����)���g�|�ѣ��T���+b��/�(��ߣ�\H�É3L�p��w)�Y�9K�{:������ޫ��_��e3�Nܭ�ܮ��"G����<ώ�_
���J��{tzoً2���`�ɨW!�S�e�%�v�K��*�񬥯]=�u拷ga�ͽ��8�*�SH7j�6�Ɨ9��[l6R�2F�Q��%
J�}Dv�
��a]���{�]��(��h(.`KRZ휮�P�� ����G&�ꮲ$��áX�n��w�կ�J낸���4�և��ь(�Mm�5R�`0�������F=��yѦ-*�}�qO��L�Gâ��ZA�[�9m�\t�+����)$A���K�;�R�e6�jc��lT]����4t�څL��Gv,��q�g4����y�ho�P���0X6PY���yk�� ��Yt�ںu�z9B��;�t�z���󮌥2�Dv�u�ٲ�j�h(?)JP�q)iF�e��yi/^�7���޵.��vs��BB�S�����h���),X�ǹ������*n5/s�#Bp��+�|+	1�F)�I�<��R�R��$]���x����I�z�%�^��6��D�/��X�clNS��
ڎ������m���X4��4�E���'uf�!39A�&��uHN�u��E�իd�O:��8u��>��W����x��<�.u�\�BCCv��l�y�:=��k��sw���
���[O`ʷ�a�ܖ��բ�u=Sy�w#�o�:䛁�Y�W�\[u��ɚ���x�z|��hɷ����3����2N6�{��6���Z�}�1x���Ұ��٣];��MvM8ڃMF��1�-�agb��b
'�H��.7��:̽pn��U��9�)(��9*�[���Zv�ɝ*��cu��G��W692ѿ?r��_iI�[�H��Z�ٚҰ��g^f�fl'�(X@ꉲs_"���e��p�BO��Y��^U�b����3���������z�r1�SE0oU�7�����W��wةe�7�kߨ�n�k�Ï'��b��O򋮂��yPZ�ޡGeU�ѥJu��]�*۱$7��\�,��G��]�6i�P���`�떂'��%���Ǫb��H��ZDpʥ'h���:��uH�i���m�qT��
[.�BB��Ha	A�8���_q��b����P����BZr���N1kT�����c��+CPFѭZ�ǝ.�9C��)��瘪f�kN��1�5W[�gA8�ټ(<�Ae.�h��m�ۇF����ڥ�sPcXu'W�s1XwvF�iơ��7�Q�v�
�Ʈٻ��Rvv��Ϫ�>��5�գY��g���z�f��8$�{7(�ݽ�׭Q�
h3&<�C|RD��"|��!PkN�����uB�b6v�Uq�?��_Vʰ�۝@�968��mZ�Pk6f�1��T��g�/<���>�o�S5��]�� c}8���&�l��Iˉ-�$�m�}��v�@g�0� wc�_x�ӹ
oX��z��szpI ��2���/6y��ew��Ÿ���>����	����9��|�r"3�|P�}j�!3�\.E:��W��u��5A�{�Y��!~�5/��,�������J��3+6���U��;�]�u��\T�#�<�V2o�g�����[�Q}�}ٝ2����c;�*WM��������}%�>� �O[�܃� V=�j1�يM�u6���n&-��.$!c�&V�!c1�4�mh�	(��r^�B��־��O�͜��k�Z�!��"	�ͮ+���u�y�d�3�;of=x����]U���ZVfk��ٱ��s&��۱'i�v͢�ģ����O�
��� �_�z�X�03ν�9�E@�û�	��Z�����w%�4ц�lb��E�nj�S�S��N&

�Mr+�el���xv��]٪�ۊJ^g �vp �|������<���� p�d5�6�<�]W`�d��b�㲛�-�`�u��Dp�u$�.�F�
���pM��TX^��������([I�#i��	ta]��X0��ihKP֎볫��hѵ��k�Zph�q�{����F�zE�(�AHH18t�X�#ln�ANqy��p�|'��u�������8�q,-z�7�T��P��)�묮�j��`��J��i���J�h��e���۝�^s
 IUM
�g�Z������n
Ö[�HċNͺW�4|�g,�馯�oW�6�z�{���㬿7E�Y��F��GvbCM�=�"f�N�ʬ����3`�X���a%��;�޷���<��k^.�ٚ.�\h��W:��Dv��;GL�饘�qy�m��+^J�{��X�οq�mK��%|ϱbAA0�P�B�EMU͝s��
N[��I�D{6�*a��S2@�N$���R}�J]�r�vkP���1V*Aqsb�m�gSFL[��=!�a��p�
��(뺍���ј泵n�g���]<ţt�:Q�i4�}Χ���}/���i��C���,j���^w�jH"����O�Xz��o���el����|��T�D:(P2���M?X��A�u�H�2Lj]]X��̉!#IF\f,ީ]\�xf1nw0���<ZM�}C>�@�]�*7��d����B�iK�N��b�	���.i[���/_`�0�˱n��<������n��,NS�������.�<�ؔt����\���F�����ӟݕ���r�9x��k{�;�Ҝ�V	��F�[�G��5M�����#�g6qtY�N6U<s�8J�����B�����t�7�k�=:{|I(��a�޽}���KX�El��r����HY�;,� �M�awe�{.�姈�&��w��������Uu�3��ub�ꢭ����"�f��em�`����-g�۾1x�qC᭘��S�d���4�@�gP�Un��#��h�Œ�뤚��dWe�g#KF��RF�e|�n�k;�Ƀ�;"Nƺ�f�I����Q�/fY�d��Ik.Ԓ5��{,�b���t��0u���6�˧/ua��Г���V쌮yB����=R�tx�Ϳ�k}n�-�b��@^�g]��ȗ�P;6�ǭ$�@K�KoKӝ����׫N�iqH&����Ӯ�S���Q5FbxCZl�R4[f����JJ�=���!l-iP���j��q��-�j����	�&��k��s[V�˰lڹ��2����e��`�1+����K5��Ĳ��֭�]n��SQ[���=�I7'E'	��,#�ОP�l-�A4Y��s�ܐ����+y��dd༺�$�C3G������t�܎��;%�j ��s�c0ONtf�ڸ�����
��@r���$t�C�	���&j��:2��u�HB��u�} "�'P��AenM��}^sG���G�g?�:Mph�H膘L��5��H�T��l�yL�ł�O�+0��n$���Q1N���*M���!2�0)q��,\����:vӰֹ�k�'U��ퟏX�4F����5zLg�x^lx��wX3�`N�Ё�݄سJ����S1!�`�A���8�hwu�vI�ۈZ�;W�V;�S��.���\��#�ia���꾨_pCn[V��m �n��� �ԳZuV���dn��f6�D�I���=��+�QT�$�k;�v��o��-�H��kOv���s�==eƔ�O��Fe[4�y�GV�ӄ2��dY-�
��"�d��c�H)6*��Ɗ���K�@���{�1�41W�\�k��ͧ޼ ��_����A��H�q}:S1��������@�g7Z����jc�%r�ι�YE��K��ޠ >81a^�aO��+vWi�\sH2��wm߈.Y!�	�A�-�d����̷>�g웁	��{�oW�:�߱��/� Kl�����B���^ܺ�S$M-�tN$�U��	���ǽ���<��G����zV�XǹڈI�Ӎ&f�yLWen��������w�����G�]-��Z��Xv�%rR�'�I\��C��:���`*T�?��5eVF�L�;3���M��F�ܶ�j�`��J��%��e�a�4�N6u=ݛ���)n&U���+�2ZZ�8bۘ@�Wv�82#�O�. �g��ۡ�h���#L�wC1��K_�z8�O�A��$����
�::�^�ȶ����(���j����S`�ƒ�5��rȬ�^H���)��!�fF��+��qۭ�Fc��*yIQ�n6�l�
����H��z���!מ-V�����x�"���"��7��0��ŧT�dZ|�����S!���r�)ĳ�({�z�\:��Y��f�k�W|�eP����BF�9����\׷L�]��&ɩsh'����-�(�JH�N��z���c/EB�QWg���f�j�Jn�F�O�1��ý-6���?0�Nm�ɧ]&�j�nΜ�$t��iJ�ɦ�yxy�[��i7�h��AF���PF�Gm��Ȓ!�ZB�R����������b���y&{�qN�a�ϱ�n͎*�i:�rF��w�=qT�!t�]_N�:��L����ָ����1@xq��E�*0� ݋��X�}p�H��"</
�M�/-��S]�z��;����s�����-݇B�i	�q*�j�ߗz�*Ț7��}����/��e;4?ޟ��xmc=º�h�#N�#��2TW��L���v��Cq[�;�<1��XgH>����	�.�=��Z"�$u�aZ��7�p�wrj�vW^_ �Y彨�,P��Q|���M��[���B%$ ���8���W�em73�\�,J��G#��P�v��B��e�i]'QZ���<� �F�w;��w,��%���I�H�g���kI�^��X�U�wR����V��� 9��rfo�R��⫥�Ћ;�y[ѷ����+���%�W����'O.���%�{��*��Յ�V1U�̥r�WV���e͞���Gw9�Ɨ˻�r��w]�v��S�	c��3�u�`DX�w��Nv���]GNK�y��/hZz�?!�LSy�l��un\��݉�1� 5��3���Դ�����O)�L�����|}���{}�_�         e�   �k������,�0���^u�J�kG�Z��i2�]5fJ��ݝ,�3Z.�/Y�h�ĶbVX�T���o%fP-��\9lCWL�6�4�����:m[j�m�{m�kU��s���G�1�O,���hې�j�s/MF')�o0f�����<�3�f���mv�Q���1���۰LZ;(�Rʩ���6�c;f��*�2��ڒ��l��b�j�Mk��Uh�6��T�a;��-����م��VBT&Z��k6������X+�)���v-��3-��!n�10lٜZ��4Ba���%ȬٵҢ�^G͌K������1b�0��#�q�W
 Ō�m�Y��Rg��C8�fWvM�j\v�
�ͪ#J��՚��cL^h��u�]�ݍ,-�#lEa�̮���sz��7k����-��ʕ0�&��,kc��ֺ�T �ձ��a�����f�Λ�[\Z�Z495�D�5aM�Uu�ܬ+]#1��·W��Kbj��˨R�l#�Z��gG]vss�^��	��V���b�q#A�(F�LA����s���O��w�.5�5�t�Z��[��.��M�K�1[[�+I@�f�]s��qD�2���]�`d Mz�ЍB�e���:��tηWq�\�n��P� ��f��X��C#ulԙ��Ʊ�	ť��8꺙R�4 ��8pg�%�3�`�e�Ֆ]�1������yN������8d�w��7��^7�F�K�l�[�%1u������60	�C����k��pY�#���"��e����Dd,�aB�{`ǵ��뜽̒g=���-scfk���\��2q�9[k!r���E���7��G�n���v�\�Ȫ��%B�)]x�v�q��,w<���{�cM��ե���2�u����?M��Ky��f<�o���
n۹۴R0�a��2}�K�ݵu��"mg�:�V[8̄�;�2빚�q$QV�I�ݕ�B�
�b~�Y���o=��v$k���㍖�L�;�ZG��R{���r�e;r�KW���k:��o����3x�SNIїm�����H�vv�.���,[X��DA ��wQF}��KP��6���[�19�d���r�R6{*NY�0�G0G%��M�_ ډ����JV$ʋ-���Y(E��<�z��vMB�e�70��v�)�K������V�-2�R{�"��>[�8��5��L�6�^�˝��ms�k��J�.��N��w�G[X�����"6�pɧ��q�:�TUmCM�u,���/�O2\f��{iWq��n�ޱsB'z7+,��Ȑ�j�WT�	�I��m����䶣�\lU=�~�-�*��u*����o���xm�!_s������>�7&38{���8��*5�L��Y=�ݖ��_Uo�xA���uw*��P&5�'��:M�|��<�zg������q���Ӊ�͞��W�����&V{�-��k9:t�*��WF����b�x�K2;E�w6�-֛Tt7��F	�F8��U�Z��۬7�J�j���n�	���Un�,��-����[�qBp�+��~c��SP\��J_]�מ��[��_��c
�z���S��P���w�H�*[���Z��Po�E�!Eq��	4ӑû�X2b�wڗ�����3=v�%k���Qn�n���=H�*���X)|B�ڽ<�ڑO�*�y�_o��Mev#.�E�9���/pI��7#��G�3dbV�5���}���=����0��i�3�(��-�AGm��q�ce���_a�˺�z�cvB�4��u;�dΒ�	*�,M�c{����)fHsӭ8�_�Uj��T����)Ӎ���U��ت�h=꘩5r�����0�i	��Vv�������$,����q�o���uI����^��u�{���r��`�z��z����<	��H��&&{����\�=
� S���M�%�@fO���*�pX��q"Q����#-�wN]wb�.�4�.��i}��38N��D�����<��9{cj���3p�Pv'���^Z�s�+}5�hO\�:#<���?@ �	y��id�:ַ�C4��cA��k���+�At	�h;�%]��R��b�F�-��¶�ٰ��U��tu*����uژ��jԺ`�f[����`����zgnD6�6�1�w��/X�׋V:i�|�M0=�^���q�6��k��aKi��[�Kh��?����^~c<����tJ.��rb�xӻx��Q49L2�Qa���ǽ�M��f��rg�g�+�#�Љ�W��IP9m���{� ���Jl�Ӻ�c5�7���.����)T����t��c3y�L$�}
�7�I�
i��A0�鎵͡�����<E#4�y��܈�s
�k	$P}�{P�aa�v���E����g���1V�e_8���l<�s���*�D��/�U����4�%���- (�"�ƜIϥn���8��sn���lnM0��"#~C-�ۺD�j0�k鷆�U��ZγN�l���Y��s(S�5�I������u�5C���Z�=\�<�G��:��)]k�XH娢҈!w�s)�ᦺ���&H�e���j��(A�b�X�YSuh+����܃��DK<����:+�-��Svm�@����õ�le�=��iS�t5�}�o��j�0Z�}1G��t��%>1�m�;֏{�iW��΢����j��Laab�>��h�yS�q�Іc�[P"�)>�C	+D�%�7Y���f���6Fw
�S�<����9A5�'�ݫA�t8�%t1���4��j�,��9^�J
���v��̤��x"q{Еz{"�C1�b�2����B�7���KXm�����8t���w~��S��=� ?2�1�u��f�7��oY�+���]�;<)}���R��OƆ�)p�%�K5 �\��Z|��k��X��Y�V�ǫ.�e��.p�7��*4�����xn��WӾ�0m�B}��q��.\8�"=��,�Пu�ޡw�B��������i�K�n���i�1Z��k��^%���@�mZFo?.�C9�*!	
I�9"	���d�iN#=QN��t-6����79�QfqU.Z�6<H���iy�.<[K�N����p�h`da�;�wYE[v`��S�ڵs7�Q��1��"!�(���HH�������E�
�4^2:u�yll���&3�!K��Ȗ��1�;�ٹ޷�k��4����)ې_I��K5.�x-�4�V��F́&,����G]���	Ue7 ��i��C��-K��B�ͽ��v	KP��%2	�q�@���1wf䅳187�Q�䙣�>�'E����|Yx	��_%a:�5�ợ5���D������0��wy�(�j���i���O�3z��JZ�$䓭t���$��FR���"�%:��a���b�$�d ���o��\P�"�3s�z�zŏ�I\5����s��>�n��F# ����,H/���(B4���.����p�[����5	?^��Ө�X_�պ�y��L��Ǎn�A�h�/qfz�W>ۊ�a=ݎ�'�D�[�w�I$�HS�W�F���u�YjA��Xe������fiTČ�kt��ή�,"l]�l�3Y�^�"�������x��Qr�H��c���Uu����u��r�=�zn�O^���fXr�2T������|���u�$#�W(�i#�nv]R��6f{���~��F̏&�C1��7�rs�kzs�����$������M*X{d;�x���sA��Q�F:�Wy[*��0�6-ڡ�m�a s�1�Ъ%H�m�Fc8�"����;kQa�ͣ�=�-tq��"�[�m@`)W+6���s>�W�;�ᗒ�����1\��b�	7�	��I2`0Q�n,cX�TI��\����]BC�ż�ٽn	�9a���b����-�b[�lFe����K6.�̴����݇w�ޛO/P���lbD߶���5p�zRR?͎�E�T4�G��U@��ܳD�2p�)Lp��Vyc�<�^���c�����fe�{�g^:�k���_N�
e��:D=J��OE�J8㋵#zܢ#fAW+(M�Ҿ���;G7B���j��+�Ȝq��]��'7��C��Dl�IK6�tK�<7E���i圻7�`��:�DbژI3N��م �l�O���li��3DA�4�嗙��2yd�7�GE ؍�!��&�,!sR��D���MYUn�g�f�ͻ�<�0�LD�Нm+�ŐV���
�b��Ю�;�3j��B2v'��3��7.�@X �}3-��S0�ҕtS?:�r�)�-RMG��U�Z�M�ܾ=S~�+��>��9�X�<�M��hʵ��hrWխ�c&'��&���c�N::{r�>�̶%�+F�j�3����y1"���G:�j�V��]Yr���Z��|�X���p/uk��.�\��.��>^��qy-{f��W�<�t��s�R����R���h����4s�9p8��v�E�C��
��1l��R��7d^�"CC
��dkW�zm�Yo>��c"��F�:�?�_CG�W_([�+�C��՝�âzC�s���8�)W���u	q>yeٛ;��E"�װ���%7ޘE��y헍J���\�cz��k����o^:=�I�kc�<GiIl��r�I�·r���$L���+B�|����+�w��8#|���Aл']����nwKn]go��)�j��:��{/V=w�ѹ�-��:���ʸ4h���:x׮î�]����k�h5 �*#���j���5$B�-𲮊1�x3*c���Gǥ�Nil�����n-Q0Bo\�x�V�y���g#����
*�g�VJ��}�p����vU�]�:�Y���4�o"�Ymw9O^���'ϡ���,���  \�Ɍ���oˎ���CK-p��
�lܽ���nà���Z�Uؐ,Z%i�$A�TE��i!-�:�,+��m!aR�7b!��wAb�k�b�	��p�%�x���2���5֒a@�LQ�]:[ܩ����[f��Ĭ�i�����>���{<o�r��Xu��Խ9��GF�^�z
�a�ZG.(o �N�/E%��r��;X=�73z,��}�J�Q�[ys4�.��wy��b�:��l�fwk��X��6�E�Ĥ�$%H@B�D���S��L�������g����&r�K�䎅Eu]u1�BP�HF�a&��0��Y�K�%e
��[�|������Fy�`�Q�/�(���]!b�b=.ʸS���$�Fܔ(d@芠Ƴ�K���؆$J��w�I�x�q�����F���c��|�<��b�N��H�N���^�� b�WU�yL:�"(��\�)icc��TY�C��;t�W�6e�a��8��w��¦=k�{��=n���u~�I$�I u$�4e��t��6�[���Ve[��0����M{ ;#,������Kn؆���sVe8�Z�+CKu�F�fRb��%�rYdcz7�z[!�^jVC6[�B/4�/�E�n�������n�-�.3�F�-��e�j���5�o��I�$I]j�R�r���51��T�PLUr�n�7�IM�.D�oϑ���O���>�'�L�Y����[�sL�LhKL�.x��!�쮼��F���,�28^p�h�# J�LC��Ɣ��`}Zح�i$�V�5Z�%�;kL	U�&ʺ�0�h< �G�����~��ן$ �;5[�]�\	���}ݻ�Y~9#��HWv�'�<C�
,5t�����Fۜ���tŦ⤘r~�U"�����m�wc�^K�$n �+�h��ƺ>6�r�]#���T��\9h4;�F���6a=ݒuV�Q*���dqל(�G��]�=�5F�̽�L��s;h�>����"��in�J��8;~�T�c�c����V�t���K[�GG, ��&�=�ED�Ř�>��7o4�Er�=�R.�j%K];/,�6^ߍ�wu<̇t&.�/��v��g\��5�pI�3�v-8�A��%��l��^�&��'38nvLY�]��"�l�ϩ
ׁu/�l.F�&Rd�� iB9�Zh;Ic���tң�6V^3Z�c{��Q��S���]�ջui�Y�v;[O�&|�r
9Jh��}�aaU"d|e��Y]�A�����y��:;$�z��-�Q���=�Dj� ����2V��]:5{T��kg�8�ۦ�ҭ���+"�xK�e��\�K�.P���S�17����މ"��/`�&^�v�ΰ����[�m�^�.kTÛ)%i.��V����7|���Y��˔tg9��G��v�5�R͎ߟ��~��!v������J�ҙ�J�����iF���m��u(r�������X�c��#�<cC���;Iۋt p�n��{�:u�JT�K0�:��ÝJ7j���跹əݡ�b5D6ԕ8�Yϖ��U�� ���L�L�|_2��u�R+V�?Q��O}�xP����tM�vHv�
7b9����\)�ׁz�M>�Ԃ��V���ųa�i�\D3Mo#�ꤕcR�
�J��ϡ��,vP˧�Y�RT���k��"qG��)+c��"aD([mdv�2��6�kc�XS^�Ȝd(�E+�I�ݮ��r(>��-«�}�G�vkU��v�ѕ��ch,��R��o6o��Z^[��M#��So<�[�=��_B<�-�'H�R'шDVNN�5y]%�\��!b�3v�[{�+����k�T6����*���S8�:��9��G������� ���јZ���s��=��hQ�4�D��^	��N�����S0�Y�.f� ��Tcj��/��� I�-�-]�/�_;�	�=7�O7�Jg8ܥc���U�������[��Wk��'ky[tY�m=xA3��;�RE��M0��@`�-3X�m	i &K��A�jVf���Z0�.��0Ѷ��Ιn������/I'LE�nI�CK-n
Mi�g�5�ķ��%t�l�`*����aWj�TK%���u�%9{b���z�U�I�[m��h�U/Rw����f��>L�]��@bZ�8ŕή���Ӡ����$�j��)�)V@c2�U^_����H r9n�7����)�^-@�y}�7:<���Uw�rvp-�Iȣr���Kd~����7�
�1��rͧO�s�k7�acgAg��/	��8Ӭ���[�հ��#�gL'o7�r���k��w����X yN�Q�"٦4�qQ��r)'
l�.��9��n��u��c5lcB��P����9Hf��Ͻ y���z�	u����O�1�֪������WW3���7��a�M\����r�6�{
��+���U�wH���������.� �[E���kP�ʆL�)|�
e���L�V�nT�g��^�f�֔(]�.�WG$H�T���U:G�˸�
Q�J4!�e��4�<���r܏T6�C�i�a�&u3�0��K��#?[\_B�|(��$Z�kmŒt��&�|���$F]�v�-$IS%�Z�A�mmڳH$���{�̔"X�t,z:_�Lm�����If�w���T�G5�c0��9�+����B|h�eV�QG�sU��n�v��c���8U3���UZ.�7�.C��_h庰���CD�s�I��#D1Xj�ә�3�9�am�װ�fU�'���T)Z+rJ�hAD�;E��2k:B�7rMõnI7��43E��K�Tt�$��v�V��vN7ۦ�y��&B&��lQ��(Vk��ɤ􏻉��VlF�1@��$��)ud:'Mǵ�8�z\�j$����z�x�P�[O3��Y�J��i�^��7|+�����w�ͮ�# ��ҹ �	����+�)�̎E�C�W=����d�l4��9.Y�$���ҙ�m�̫�8=�+4,����l'��]��'�5z[��\+k�V�GT�4�I��+��0�O�	2W6Y;�2�ZOI�n�`�o��Uw}��lY��D�в��u���s�X�ЬAN4`�M�F�wK���*���QQ4�Am�8�N��]g�R��tQ���B\�`�FZ�l����Sʐ��cT��.�M��vd��<�y�Ĭ�k�1)�
�,n��D�R�;Ǹ�&V���uӾ}v `�d؁�Sp��p����p�L�}j2��F�UP��8�n���������^��h�F��)�J���:�^��*�_�eL�;�`�tb�,=�pψ��A2e���D�T�qJk�T����Ԙ�e$+o�-�q�ޣ�`{C��O#� � Q�(>B/���	����Α  �   I$$�4�*�Z	C�C�
�}f��B�[�)L@�|��	̸���@D"��A2cc�74�SI���F�ED�l<\��[0b0"K11v�X�"7J�9���)�B�㖏�Xm6�3X�oL)��nT�ޅoB��D� ��.q��ؚ�R�5���"�� ��EU(�"���� �E[EDdDB�(@-�d� 7 ���"���(#b ���h�%(��+���h�V@��@IhQƥ�1��7��y��p��[[W�oM5�sG2ױS�QĪo�b@ �%%S*(I�B.�@Q`0�"���K$�e�e��hH��H���& )��R�o$�IIP��N��}%�d  0 VA$��mTU6���/�*o��~\�D�-�0�)dC�N�`�]4$O����gPZ����?�q���?s��A�)���Qb��X��oP�7O��K<�J`�?�!�����Y=��M#�%P�Kw�����y[�l�.;��`"4+HnPtNcd�*�]�;���	@�D
)�к�C���	r�'1�%́qw˅�vCи\x��q۠l�lC�\]�Tg�zwm����<�ܝL>��$C�
v��>�c�F� j��P�� !�-X�dW�AT
_�B��`�@�Oj���S�O#��~A���<�����&�s)<Cu�A�=ޑ0п��+XC>�́,.V�)|��=~"l��.��� d�NHt�H��0�RE��|���ʈ���`\D��.BI'��}X�=�Ct>_�s�KG���X�����p� �n#�����{"��z��-�!B|ś���ְ��XVt.Z	rHB���,E�	z��J�B���i���C*����{��q�j�˛BR��Š���,�������T���%��!�A� HH!�+Ĺ������l���LzSb [F?z���4[���>NJ(�h�%)V]	BR��ȸ	`�F��R�IjJs���"�H
�#�
6mq, ��PY"B���4Ţ$#)�JDK�7-�D�� F$VAD�Y P��N����\[X\�|���5���?�8:\����u�����LO�Ȅd����@��@�����FnB�$�~�������Jw�kEO`�=Ȫ"�)���d��=�/����T��p~�"�����GX��d��KC�,'�����t��{����`B	O�	@��ɰk�p:_���X�nw��">� �����D��(��%%���@|�e��H$ % 
���i� zB	�A�Ji"�৩���	�t���.�Ǜ�2|	P�/����F ������_!�X��s/`��B!��J864"u�e��O�`�A=��e;�M��XO�!}шA>"u!6;�w	� ��~'�N�I�g�C�|���`�ǂ!�`v�@����o� ��9 B���*� �:�@\EO01�0Q������Sҩ�K��.9���ؽ��b����4�����t@�1Vϰ|�B��H$P�a!�d�PP"�r�*��'�O��������w�F�� $=i�!�И�p!b���n���1�NGh	�����%(���r(��B  ��"<D���Q;	hJ��R(�d`�	��a�����ȑ� ��J h�'Y�g�&��EU0�E|�|Q�C ]�;�nX��� �}�nn1]�`�.��0&��H,�?;RH�B�-T�j��	�PU�B��@t�./Y|���&M�[�l�p#B�cp.R!�h�d��	��\���\�� �܈��*����A���	:0n�r� �*�k� BB�R/o�L���/W~A�.	�p}a�@0�Y�!�lE$Q��Q@�����,���~�;����C�=ɢ ��<���ǽ���9;�@ޖ�k����&�~�4�6a<K�����[����q��!~�Q8�=��$�ZNG������ ����B'�D����_Y�"Ddns����&P�9���7W�^��N��E�T2�=o�֞�$$$$!A%Ҫ��2D�b��*P����1j8 >�DU�� ~�}L��� �9�����$o��PX���/Py�kT�b�u���&	b���aHeA��|ˈ���_0d�7�x`�r������HA�KX����Ȗr{CmL;k4��"�w�\��F�?TG4�����{'_�!��w��@�Uϴӯw���|�	���, h[�1�ht=28	C�Q@n�^5�8\K�)�Hp�6�4rSA�$�@�I%�x�;vz�ݝ�ƈ�|No1DU��?4r�\���y��*�V� [a�l@9x �	��sA�.&��%[�j��pdM�� �>!�Se�6���l�_�jN�yBZD�"Z	"�H#g�((��/'�&�{zD�&�Jr2#�_p��tr9�8[.	��Ӑ��� :�����y��z"�@ ?R� P=�rW�p^��'�_�v4�h�KU�#�;�~��u�稳����� ���Ԁc�M��,%�����%�,9�&����9%���7��G�$�zg%~0���r=��U�?Qp%�$D�=��VDn0~���V	Xz�<�����O���ܑN$,"U��