BZh91AY&SY��E�߀ryg������?���ah� p                    >            �          ���{b��'��%sj�T��P��^f�
(��y� ]<� �9PUݹ%�(N�q�*��T$*���G\MUU,���݅
�눻j]`%��vVصqл����.f+7wvF�97`h[�4t�&� ��    �ht�95um ��`� s@4:j��c�ҨlP�4�2� n��ӪP\����ri�)���ih(�F ]�Iv5�t�+��ˤJ�*�5NM �v(���WT�;:٢�5@ݸA�ڀ�j�4BT�    :�4rкԒ�j�+CJ*�6��]��l�(e��kY�kfT�
�V��;����EjP���ҕM 5�&��R�V��*�ݚ���
�A0    1��ݹ	r�2�X�N��$�a5*�g�������%EB�m۷Tp1kR���;�R�&��I���wu �Q�J����    ��)+MA-�T�F
0�t��n�UtS��0RF]rىU�R�Ui�,�T�)*�Ȇ�*�k�À@
aD�H�MA3/ =        ��T�I�  A�h  S�"R�(�`F   4�2dшbi���4�&&�h �?&��I)@4   h   "L��M4�2C��6Se?I���OD!)QF���1 ɠF@�M4ӻ�y�)<�>L�z�5{m1+|d��s����d�qx2�=Ȫ���G 
�ࢨ z�*m�����FTY�!A�=���'�۫����lz=Z�:���������;���,?�|�:�D�BA ������� ��.��#���Ŧ�A�u������t� � �@@ꍱN�%D>���ϗ�g�������'��q���3���~_�?t���;�Ds5 DC�U_N�h�w��b���6�f�>OEy���Z���#"Up|߳j����ێ;;~�^o�mH����%i	#����,���7�e���=1ܺ�0ek�6]�;lX�M��7�����	8�������\7A0f�	,���
ջ9dhn����W\ �e;w)cL��9tJm���v��g�'v�չ֬%耓�,[Won���i�Dw�!���n�N˨A�e��DD;�U|n�y�sy�)R8�(���}�j��Wy������Z1��f��S&�7�v�b�{Z�7;�����Nk[�s�{q0��+[����Q�̎���j�ۏ���޶�4�{+���nZ�6wspo"��8b��p��|�Ɗ��t�|�s�Ѹ9��[z7#�ѐ�����5���M�o
�v��`���w*��٢�W7���j�\<syeh�:���"a�+ӹ�n��bˢ����Ś�M 0�Sቖ��hǘ��j �y�ܫs�.o5�sXk�؝
0�Y��;݉b�2o-nJq��7v��{j�Vo9��ߵ O��K}�** ��rt��a�.�6����co �寓\��Y�܄N]Z�`���z�K�:pN��W�V�{W�t�h#�vl�b�a���\������,7^n0ӮԬ����M��}���2�R�1������{dRl���~��e[BA���	+���+yS��t���"rʔN�N�F�@v�n?�X%�x�Cnj[�h��(�F���7��Xݱ�=���ɚ�Jc�^�u�&�]�r��W��zѻr
��v���:�#C����Y	�7pJ�&��ı���l;fo=!v���1B���5���M:P:�i�ܱ��œ�7x`��y.����2��v�aۛ�y��� �ӊ�_^Y�=��;&��P�[c~9�nK��N��+sQ�Uƅ	<��㕒���\��v�u�o^c�(�%�g�E��`�<Sr�p�םxu'�d�8�LۣS���[)
�S��#��Gr���n�S5�C�^�$����V�����~+cJy�d�s�����9�*sP;��=;�9z�d͏��-xB�n����P����.�Ҿ6^�wh���^]GPaogsƦ��od�]�#�6O�w5��co��2ov��8V�ozk0rm�s
�{
�ه��Dܥ׏Z���٣Z��f囝�`�a6���Jf#���ȁ3n橝#!������~$�3a��^(Ѐ�%�����+z�Đ[�ᨊ5���H�+E��;dÝ��~aө��zC�{��-�,x�(x�:G��8�Ҵ���Kp��u�6M�(�݄�o	@�+����FIPR͸�}~�E��F�gb��Y#�w!�������ى"6!�c�.��O@�^t'��2/���p:�#װ��+����4���ⷘ�G�5�m�����D�[9��W���\���H��]{CUd�[r�L�f�v:�`+v����{h�Fv`ՏN��0�|S4�� ފ��֢Q�Um��:mf�8r�v��p�J�r�>��c�#��%H��p]$�-�MaU�q��Y�u����.��J�\ �wx-�~���
����R���b���3�c�c;n�����
Ѯ��2d�JLHΌ���
�"Ό��U*9ro�51�+m�{�������ܛS��v.�հ!+�iD�7�<�@r�ɴ�rB�w���-��P�(���/�'7���r�<�KR��z�真cs;��F1[�$wM섀ܨݙ���K��N��f���Y��9d�W����+w�S����3�����p��c�:H�ݺ��7�Na��$&�Whi�F��v7;�)���V��9�I�7�������: sx1E�Ʌ��[V�V�z�홪)���֧��g�+rqsfol���h�"�8l�wэ��d죵�o����u5�(wn]��c�z"0]�t�3u$�;\Z�p�(�a�R,N�qY��j�f������%8��;^�u��n��ݶ\�4�A�-���^_.�J�T3�
� *���ز}�~�ځ��;%}��!CGoaZ���U�2r|fv>zq6F3��ʖjם:�;u��K�܃U:�#T��S_�$��*f
��@��"�����A�7C��e<��-@�uo@�n�c�\�B��9^����fs��M1О8�}��7^B ��݉�߫0:f<��(0�c|��qǙ��nj� �s��n¯W�N۹6��,��f�ͺ��Nt�b�㯴��f��~�1b�y�X�&_q��#I�9!����m���;ƏQ҄3Gf�1D�i�s��#�b�#�,B@l �3Q˪�((�77��X�ƤK42��%�<Հ���v8�s5���]�I���rŶQ����n'Vq\Y�ם;t�Ѓ$�	g7�Z�e/��ě�ԵiR���(���#�A��W�)�$�PvW˕�3�nNͣ�%�����9&�̲#��P^΅H�{ᒽ1��wY�t��^��\���2����e�ɢ�tn݊�Iى�9�4�����h�,9�&���Y/ �"�[�j�u	y�É�D�o�gC�s!9�3$�N���F��@�YV���M�gw�.ʖ�����Li[���6ps'��]�yؠ��f@G�S�Y4�Q�u}D\�Ap7���Hʭ��-�2�;x�Z;�.���y3e�}H�ͮC��u%'�Γ�K:{vL�o�r))T���:���@��"�5a�mڞ,e�{7yoj�����*�k�^	1�E1�� �'<-W�v�N������2��P6S�B^و�o�p!��֣�@s�o�]�ۼF54jE��XW.'RSQG��y����p�J7{��Y+6mˏ����
+�
ͭ"��y���Xw8��G`ޯzf>�I����r�^SxEf�n�)�w�ǜ_.�F�F���_M�Zv�N+�-P�K�����e���a�6��a��3�ٷ(%��\���}��]�,u�I�6hY�w�:
:{��M�b��4�p�e��B80�W[�G���|(ÖB�� �euSc�X��Emڷ0r���m�;����h��g7Y����mc��&̶d����F��n�ݸ���Ȗ�� ��m��L1�"��~ gj�l��m%�l㈾h�s�\��\�8ě�pkA}�诞�a�����ȏ�M,�9�N<��Mvnh������SUѩ��cѹ,�X�@v���u�I1�	�&�2�y��b8��B�!�a��&����\'����9㋲�gs
-���1-կ#��$���Cj�d����2y�����$ۨŠ����\�51ŋ��g1a�*���w9EV����ۺ�E�l��/�2.8t=����i4��ɗ����`�^-K�����1�s׻c�Tȸ��8r$�5�z�]Wy]�q��K3A�L�$�)�V�Amc"���X@`�U��v�$�ővޟ\�u�����P�o=)��b�pn����v�8&�ܘ�xro ���DR'�2M�]"� L�E���GQ^n�'��1�%�Y+���5H�h�i�H�wиγ�;�^�2��7�U1���E�<y@y��
��콽׸v�]�HM�>>����t�k#��-�_+�u���sny<ܼ�l�����W�: ����C�_����L
*|W^[L]�'�R�n���<�vLu���gf3�g�ijY�iE�����h��5��Lm�b����������������������������������������x�ݡ���|�"n�6�;m��s��t�[�,��أ��d�3����`�Sw	���<ۗ���>"9Ɏ^��	�ய>�6r%���x<�3ۭ�ղ�۶wu�ln7g\fx����uu�Ż[�=��W�Dsq�q��ɝ�bES���M�؏����.�烶���:��q���e����Od�N�F8��s�[���x�1��ץ�Ҽ��iy;p۰�X󽽺��glu+�Mλ��iB�+���`��޳��Z�Om�nV�(���O ��z�X����x�^۷Q5c����ŀȵ8�Y���-؃6�a�Ս�'k�]=Uۙɷ:sGgQ9���<����v�N��s��zn��.��\��ܛ�u���1��]]��#���r���ۈ�Q볹w��C��w��u���Q��ٌ�]��T��m��y��ʡ۳���䚮6"���f#�3��/E�v��^���Gs�3��<���nLa���@�l����t�|�ϝ��.����dw;�4���;�i�6����v��*|L�]`7��r�� �l���\ι�-�mG=n9s��2���s�g%R���`B����&�Ǹ���=W�\v�Ӯ[����-�uůtS�O.y2�]���ܰ�+z{z�]��A�vx�Ɏ�OZs��[��W
��N{bA�[�5��p�۱�a�V��ѻb�q�t[�gGr�;)�z�nѲU̶������8]cq���2a�����TvrQ��s,�;%�۶W��=*n^�͐\p�5���:/VA睖9��κ�l��3����);Mqx�i<�"rL.=|`���� �m�qԯ�ήvgWi�1k5��O��ܱ�[n�W�e��0�����m� ًq[�F���:5�l���e��r%F��Kɽs��ܶ0\Sv��$�{<�苐����sǗ8��f�n1��
�l���훚�)cڮl�k=j6�M�uD�Sp�0[w��Ň�Y�����3F��;�m3�mӃ�tG v9�¥�=��kaf^�=u�y7�c�b׷)u����q�6�,�ke�1v�ӄ��{�+/�:�H=s�N-�wn�����{jAvŻ/���aֻZS�����݋J�v�͝ά�ey�[�;��JC���e�g�T_>u��ݡ��v9ַ<�2vMTCy�^Ļ��Q�O;�<�nv{6"�u�n�j�v�+sn�T�ݎ6N��\������`�D�vѶ�����^W�Cٓ�d���kM�\��P��=�݃�����b֯p��.�=��=�۷g�u��=�Y��4k�%\d�vj�7'
����aܵ͸��.˻�<O6ν��ݻs�@�Q��g�ζwt;v�p�烰���9��r��(�vے�'3:_W���	�噓t����ۡ�\�guc[�����,������m�=�r�x��\%��H؂�p�M�[��\p��.��C��F�ηu���`��zH�y��j�B�[��t�,n��qu���ݑ��>�M��f�]�t��E��嫛[a�9���l;�m�/�z��
Ձ����b�#�i�[������/����n�ö���L�x-���]��C�Ӗ��a�l�>�����ӳ��y�[Q�w]�nOO+�6k��V���vbug�ݮy�+��Q�&w5lm��48a�Ӯq\:�'kk0�v�f��GD���Þ�lb½U�)�[�-��ư[������Oc\� Ӣ+%K�� @��q�"v�#�^6O���vÓ��d��M/6:�л�]�)\���X]���b�f����"5u�vN;��RmOA�hظ���BI^}�[\���w=n�ʑd5�C�4�퀷96����5=r�t{��xN�������c��[�>�
t6��&��=�=��gY�l��s:('�ܱ�]�M�W��cm!���=\���Cѥ�y�D�X�g�y�s�9�A��B�\��VwJ��3�ٵ��R���dUg�np�E[k&cr���X�a�ۙ-뗛���CI�n�m�lkgq�\����n�;n�7�s8�3ˌv��kk���)�m����K��O�ŜV-��v�=�rY��c � x��F;It���Q���r�qs3�6�C�����..�u��ŵ��x�-�Jt=��۱�v�����y�x�j^��s]���x�;B��73�;;s]�ݔ�6����	u�TG%k�0ڞB$�&Ѵ���n��v1��W���<`L����b6�^��W:94�4�������h�x�8l:1Ws���2h��"36��[8�l��v3k�&�<�n���+���U��6˶�y{=��՗���x�2g���I�;I�g=���Zɐ��u�83���f��p��p�T�5ݻ[s�u��p�{]����pu�^m�ݭpq*;4�����	OPu��*���0F�<�j1<e}�>�3/=��Q�c���z���n��C�E������mɓ�=�C�g�}��n��lƽpj-��2��})��[�<gq�s�ȯ<v�XE��ݜ뎀�{I�x����Ʈ3�z��0�7Vڕ	�h��ۇ���
��]%H��8�)����"rg��{������U�oOa���Vs� ��>|E��s��Bp�<�:��9j��Q�U5{=�ۚ�7;�O+��d6��黶���v�퉞�yJ�r���\���	AG�j�z�uñ�9g�hIs��`b��w�����1�����y�o-
y��q��*�^�=�6� � x硆�� M.�o�n���Q�'�(��c��S������AT@ r�A$0O���~UG�����~�y�\L1O*����ό�۱Z�����t����
��(���1�cUUUUT=%n�c�M��Rn��;)mӹոšw��N���!�t7WL^�$��Z��lv���*u�/gk��.Z�#፻�%nz՜�TdG	��'a7N{c-��y[�gI�.���"��-7td���q���@A�p�!�޻U��9B:�^]$w�Bs���ڜu�� �L�&L�eN� �Ov�v������i��i5�Pn�;Ga�Vڮ��ny���Y����6��ʼ1ӵy㞷q�	�\T��0-�Y����;���D�������u9�z��[,p���n˺g�(v�v/W3ȭ&�A���wQj�<F�����s�Ԝ��I���r�mۭ�-�憄2����pW-<����W]��鮪�ǫ�]������n�]q���)���l&�T;t&t[;���U����Bl`��h���'5n�z0��8C�N���[T%��#)�Bl�cb�n9���v����I�1w��Ƨ���l��\��q���۳�{���[�x�gf��7gny��R���b�6(�9�dvS�i�.n�gO����ϳ��|�R��r)�圆u�=1.]X�B�/�&v�ݻT:��	�U�=�=�݊K���9-�Ϥ�x��ͬŰ�f|S��6��2�ݖ4y��c�0t�"c�Z�mn9ͷl��|��NI�fF�����w{ݛ�F�,�B���r���h��Jn�Զ0�?�[�.��N~�y[�g�o���ս�(ٿ��Q��B��2��k��x�e� !R$�c��Φ�j?�חG���-�t=V�p���k����'9�2���"k���X#�?aZG�I�y�����=��Y���+�b>�&d�3�|����Wef����G�_�/��A�{��9�x����?T�a#exR2�B҂߶��ْ/�\���Ú�ꋆ�b���|/f3���q��>ny����LT3�����H�S��b�n}�!�#y�A@���l�n�d���[y�j���-��x��:ׯƠ}��~�c`���9kJZ![G��i9ט���%e`�Ο�XU,����*��e,o��U�|��-ݡ�������j��x�[U����N�Bz1�2չ�X�,��o�<u�v?-"���6��l9gsz���ۼ�{�����ȸ�Ҿ*�xJ�{~��藄��S�����zӉpJ�X�w�K<�D�1����p����4�E���H��2�|%�j�^)����DV��t��a[���%�S��n�0��]P}ְ���L�I�R�ʠ�M-,IRJʠU�B%�x^p��:��pT�U����ڻ�gK�N�KJC�y���K�VX$m����ӈ2�%�@\@�B����&!��sOP7�XC{�c���H2�ī�cͧ�s�uK���Ұ���:~j�S<US��C�� bҪʥ
IiX��m��튒e&%�©A.���eT�{��O���Y֗�\)U�W��6���	�Q�
��-�IAu�In����UJ�	UJH-fko����?O�̛�f���B�8��hnq����n�v�J��w�{�"b)���6�ػ	Υ�b��.(j�V��\�@�uT�	��Q1��,_&���t��F�Ȅ�)�Ny����s���'P�R���@�VU3)%=�'ێ�d��� mf���DM��U[iA$Ĭ_O��t���K��s�ZR"��WZ�Dn�x�b\P� �ԉ����1 ֨P�m�Ȗ �
�vous)�J��B��\V�'��iǉR�J�5�R;��J��u����P�$B��&5�@�_s�)-P��%*	l�Oo��?&�:��\�� �M����K
Aɑ���ޚ
|6�f1��t.qn9̰v��Gh��ShN��\*��"��U��*�*��*$�@j!�y5����K.]^P3��$�x���̜�K
��K�/�cPK��1�]��<b�GJ��
���B��D�\�	���W��T�Uz�
��$�������yߋ�� ;����M�.���%W�ƽk�1���Ғ�i.���j�D6��㋫I 3�$f�H��W���T��KT�� ��Aq gyH<^��{������0�N!����6,6��!�E9�
�LT�R�%�/�7�{�d\��RX�:\stGhĈ��9�*KTڬ�0]K�#���v�J8�H��mh'M����]	pv�1Cqx����$�JC���8)+)W��iSn��OL_O�� 
Zށ9�t��s�׊���ข�.�Tu��)!����Q�2���j8�H�"�����%Dߞ`1Dx�1��.���3�Aj*f�-	0uy-$�P�TP�j���,�.b�JMR��:�X������3�&n!� GPj	�d�7\�+�%�,�: �PJ�|Q�V�T���w�d�:�P@�Z��D�1M����MD1�����s �!�<^�Q�
����p��%_�E�B b�7�T�Pm�D��!qB@�FGl�qW1E����T��;�Aw�8�x�D$�]oKd�U ���p�6ڛƋ ƹ�Mj���q*�R�j%�
�D�+*�k{���˗��kb�w�Z�m��(t§Zk��@�s��Ĕ���8�C�})�>��R�T���|��UK UH|�|�O���ުb��tT��JX&w]Un�$�cPE�S2���kF���*�RZU��UT���	`�C���K�I�n7���b�����=���c�}q��.�ma�\=n�5k�=ev[���α}����q�cT��$�f�X�	v4�}�eP*	11W�ŕA^�O��h���Wh��jH%A�����������*�K]�*��x%@�n(�v�)/�W�V$
��ȩ|%�s���FF��BU�ĸ��!A�^�(�\߸�=�Jp�t��%�*�c��U|%

����@��+^�K�j��K�iiU5�� U��w��R�|S��^���Ir��*AV-�;j�)��j�IaIX���MRҫ�1W��U��W��=��ʱUl炬#��D��%@��B�Α.pt�
�X��,(ƪ��!���f��WR@��k��qWP���&Re{|�,+;Ȭ�LI��% ���jZb	�B��9�"b%�k�U��J�if����3��$���\QU
�]�YR�Uq�Q�]�jƉ���\@��T �2�T֘��T$�h�y�Uu��u@�K�WN���4�T�i-ưT���Q�%~��-+��%�
*�~q/	 kA�>���b��u^�N��b����d�IjBi#Ğ�=��l�^�ܴ���}oϯ���M��ԭs��wU�����3̹���Z���;=	����������$�ku�gn��b�q�u����>�g vۤ�K�޻�m��u�<d|�I�'�r
��uؘ[�=��R���]���j�gzu�ѻ�Z���ĳ�J���t�-C�:@�P�&n�\Ӯ�,v��Q
ޗ��.آ���iK1�.F��ʱ�H�#{��s��VR�{�p«�\�|�J��XW
ZT֫��圷wq�)��TiIt���uϲV�Ic��S���'�۪�	b�E
�k�*�)���*��7�iZRS�H����W9�'��) �K�z�QƧ HeW�Ҿ�,��-_
��	s�r�����T��pS�p�Z}r갱(�l�H?���aT�<�=�xU�&,b�K��J�
�	�Tu.��W���]��U&7r�K���R�Ir�X�\�ҫ�ؽ�]+<׶J�����	aK�Ș���c�Wq���~�j�.j��U��1X�(w���%���菚2�]l)��I��J�J7����+3>}Z}v�D�'��:�â��I��$kH)�����#�EePi�u�\�L���~a��έ�͂A3l���:�s;�X/O�~
�c5��;�*��K1�xZ@F{�#?0�"�C��@���vy>}�7�PK��A5�at��t�ׂ^��̻�=�L�g�n�%�s�(�;|��)�_S�U��^���b���/&fmEȤ��˽�\kr�xf/O+#�?2�£b�@���r������Z\4V�hi�/���}Q~�o�,ŀ{WdxT+V�c��	v��
�K�Y{�����<F�x������!�x�o�}��#����=@Vf�DlY��.��p��{$D,�\iD�i�n�X9�*=�n��{��>x�, ��M�}�EǛ�k\ �+�|�ę^+H,�.�N=7J�|����������|��.X!�Ku�^��o�x�FB�*�G��KS�����
~����(�S���~Vj����>^�ΐ�M��+���ew8��v�cW���S��8�Ţ[HG!e��;M\}t֐�h�LK�^P�6)E�=չc�e<\4���D�`>���>�/�/93�	S��B�G;ycG=O<9�;����}�z���E��"���ñ[\l
$	�mc��۲�n�Wƛ��f�Ju9�=���Aa�+ۛ.?$lV�1������u,p�}��9=��d#϶�x&"�RM �Ql9��:��6���^̱Ƅu�y�n�������A|��Q�__��&��,�l3�;Y��:�;,r_g�S+�|�h��F�~ҝ↤����g����,1
�K<\���v���T��z1���{�
�&����͙��A -���#�~��^����޼���wQH-���unCg�\;`��"x\EB��ɳ.��ʹ�, �)��sv����6|�Hឞ��r�X��]�d��Vc���z���(�7�ޛ7��;�n:d���������;�K���b�{8w�X��Y?{�փiTG�f�a[�W�q�k�ȟ>����و���n�����
��Ӊo�=����6m9:��E啷��._l�s��7g���.GWx�/7zw/����N�U����������U�d��#���V�>U9��<�I��v--IQf��I�2�w�~�?G�������ݫ>�W7�K5^T>�|�p�Vۮ�M��@���ו����%����^6ɚ/�5�r�3�	u��,�|��k�K�JB�5}��A�-��`��I���5��!�z,�U��{<��g9;][~���/K5������#]W������A�NM1��^5���c&�7ѯ�:�\X�s:M���}{]��\b%JA���P�h�z�}l�� ۧ�&\�u����8`��B�"m��<�S�$�F�ӏŋ.�["	�{:��ou��H@i��E�j�}�xإ��9{P��`�=�BZJ�<Ŏ���l�z��PÃhnmKop���ޜ��۷�]�j�q��KhV�vvzy�����;��}�\�<Ydx�5�凒�נw X3��㓞�6��e藪��ru��q���cvV}���o8�&Zm�	�q�����ǵ��|�n�?7<.��R�M��t���/�����?��߿���>:*q��+�o�\fV'V��X��>�e�&���c�"MF�F�o%�{L�ũk�z����iod^����w�u��H�W*3��ѥ�	f�S��a~ �S������-C9!�_��L�̓�+=.OԺbÎf�<�$�"�&a)w�G��L�m.�(�y�����MA�u�1�1u]U7g��}�k_Qŋ͈�FH]c�����sϞ\έ�*y7��*����g��[,	6��;|{��������p��۳�$X�����>���7Ve������a耔B���Dۉ�?-�����S\dG�A���ϣ���(��o[}�S��*�5����[\Mx�1��q�G,���OM�ʔ_� C8��u�݅Uz��AZW��c�]a9ĩ��i6�Wx-�j�|>��N��RG<X���ڹVޤ��'ԙ�R�[2}��aB{�x�n��Ru��yų��/���yM�%Y�$�f'�0�3�j��5!j0w"쁒�^�,>������0�o40H{Gd�T��cK�s��P��Ogv�^�p�mS=�;<b�.�e�@�L���G��r�/��ΰ"��O�R\ЅEA���,�;޾��]�6�!Ʊ�b�G��ke��a�ӖV����&ƾs"C�G;r�k[�F�8���~��ҹo��B?n����3T�7;U�z�m�e�?���������\	��J�5u�^�PX��QV��oi��]wg?�{�:��哝��%�v�93�7���1<$3ݝ|�a���op-i�;�ht�˚��J��I?��b���c��D��fv��������6�=O�-�ï7n��Ξ���Ծv-C7/�n+�� ϫ�bI�ț,�VGѽՃo>8:�_e�o\w���9�������\�ˮ���^�\n�a�3<+�����+�����E7��C+l�2
��f���rbK�Ӹ�4�jk�t�3��|��O-r̓V�Z�X��,�1�H��α4nj�컃r��.l����u��k��[ル(��du	����XxJ��I%���.�
;�b�`�b��;�ټ[RWv~�����p}_Y��ͷ�}�d�� Ӱ�e���N�p�F�_��z�Kp����f�xq�&����:r��Cߪ!�Dlk���0o�e���I���.B��o�qq�U+|��h���즑��fI���Qӝ!i���R�أ�a���ā ��M�9ח�����˾V�KS�Ƌv�3"��2��ol;�{�9�خY٤ӊ�$�y;aL�@�󱲀xÞ��>s�E�T�\Cq���/����t�e`�Vl��8���>�Y�߂�{��up��*�����殆�S��=�#�i{�t�3�g�t�b�v���	v;�sj+�>���6G��h�"��@�Vn��v���Oo1۩x��.ʠ����Б��v�4bݤ�K���w�� ��s�IK��|�Q��X�jɤ-1%����눳��tv��m���⛱߇|�׾���q����������,/.Dn���N�g��	�jl�����>��Z=�l*�%�"�'�8q��A^�b�-�G�M��e�$�b� e�b��t�e��wQ��]oV�p.�^GO���Q���59�BoGڹf.	�m�`y�������(s�B���E��=Q���uC!��է�{$���k���	��c�9N��VB��:yQH���:S�e��|�	��;1�s���b�/J�^��5<C�ڣ�kD��g������*9��e/O{�W�X��:wl>�ܝo�S+]�5�F?&�xԏ��vŁl#Ϳn�E�D7�t�q�}sv�	���
f4�%Q¢d�0cDm�ܯ`�PM=��8<�A���1��W6ݞ�\a�d�CH'H��������m�b��]������SC�WZ�t\T� �Z�W�G��ګ^/�6�<�9�Tn�n�\]MT�dz�7/6v��m_��_>�K�pY���_�]�~y����d(�Q�^#h
T �Q�^G��,��e��$+8�e)w)iV!>�tҏ���%ed@�0f����/�O�N�܎�ѽ��֛�[%L��������c��K/5u�~����`4Q��0`�j
 :RZB�T��q����ܔ�
zGQEa��gIL�Q�ߖ=y��}G���x'�#
����Ae<I��F��҄LB������fD}����XV�{1b������y�ѣ��]J:@�è'u��`ۥpZ݄K\���G$*�9E���or�����rA0`�U���������7��2
p4!b�w��d4�{ίe=�x�x(��S׳9�6��+��==�܌�+̄%1�D�]xF��;TzߐD4��}�'-sU/ʈ�XQؾ�ݣt����s�?�I��O,�-đpE���~�����8#�Ch۞�4f��l�!�S��,����P��D�Zā�%{�0��ټ�",�}�e�xT��L��F���x)l��W��7/���P��A�7ں9��j�Mn�;�'o�����vq�U�l��FZ*��zE	I�W
�p2NR_j���H$�Dv�Ϸ]���A�y���a5�Hճ������k�4��N�\���Y�{h����4ū7�L�Ƈm��q��h�CCO�bg[�t4w&��O�}�G�������]H~e�O8:g[y���'sEF���sW%��$0�1?N?��\��k�v#��_P$U��ܞހze�{�wH���L�77 ���ۉN��bk�و��2�̵8�9L4���Q����o��w$��p�e i�)y\��?���#�j����G�6\�}�ڈ��#���]L�2�OȄ�`ު�Dv��y-enE�x�	S4F���Q���{D)j�:�vּ+�4QL�� �ˑ���v;k��b=Uv3�82`�in�&|�$���w�1g�)���-jm��&+����mY��H�L�݁�Ϝk���u��s��,՘�r�5 RQ���R���в4�kR#�ɚjǒs��d"W�̈́ٛ�N�5��j���'<�A�.��p\�a��黚���г�f u�^m$RĂ����iG�Aԉ��k�>�Ow���ݟ�Τ�[ ��H�g�^��ʨ%VWs;���lb,�TΘ��{O1�����#��G�ME���R�+Y�+�a��m�|��u��R䁪ղ���3Zz�涕R��B,:~�;sw�Y�:�cν���x��ZcH�g����D�A���G �.������f���f�R�Ѻ#� �jD~D�K�a��f�� ˄bDQm�;0��9��޸b�0�4�
�c��Gu��x�ˊ�ỦۦE|�`,*��&<�M�3�8|��p�q�������2e�/
-33-m�8t��;����L��Yu�|Ɨj��Ϯ�Ū�%/�,O��Ԁ��*��2 �A��9a��St�2u���%=ה�B֧�u�<ޛ�i�}������.ަO�ӓ[��cV�V-^�{�Lx����q3)��-+m�/g�L.��N�����G���XNl0���T�F?l�e̢k���m�S�Q�r>���]ض.�ݕ�<�k�+�8Uw�̆�pE"�$C,=�(㛵��d��PIϑ��������۰���S��ԑ�:�<�͞Ľ;m`���&���8�D%�pŘXB��b��u�ӸW㵰�;���փn��oU=�T4tv����vS�{p��ΰuۑ��v*���Nj��?_Jf�����ᖶ�i\�zi��-�>��k�Tϟ���>A�,�\�$Z+ٚa�6�4D"�v]�	�2E�H�=��ֿ�rKWG�&2�R��-�H��]u��sƑ�ި�.Ŧ	�γ|��R�l���>�FpA:k�ri�ٙ��=��/��c�]�]1�?\/�M�u�̋���fk�����N�O�&�#l�F���"vd��K��J���d�x����`$V��#k�=R��,�,_&ʮzpg�0=V�ts����u".q9n�|D\��kʵ�CP���v�u��v��k<k��6�xZi�����а$_2Z�͍� *�˵�j�F���y�k�����
�V�x�V��y�Y���;��m��w�y咓~�f���>�E�問���fguڱо9���yz���R�P#F&�+�� �F�V~޵���$[�\_/����A�!M����k2ݤ2��7�zX�Ŧk��4���G����a�>����m?A�w�N�����LgC�JE}f֨���p�|N4qi���t��]��*ɖN7Ѣ�uع�>���;�2 ��'*��é	��Q&��d�}@뉈o^0����%ar�s�X�d֗��S���d���A4�����(By�|�x"�w0����Rѵ�ME��1b:��9�5��v�f�M��ӫǊ c$!LC8�۵�ZT,��X�x�᳻wK_����
���N�V��A�l�y<� �u��6c�>��p<I,sy�D�o���|_6�p�   A9B�@�������=�����h3$E��\�'"�v,��&�	��;�݀kzڳ-�!����||�>�kr.�^.�(��L�^{�%��h��G9���#\�v_,{�BE{������	٦�)��8�VV�����vXw��(0��㮽�v�l�ZjgE�jq���ܱx[ǜ��\rU�v��-���"��y�B��1�3�4ε#�7d�o��Ղ��]�9o⠯�5aߖ���uYjќ�_D0�=�8��,�d�"��=������0m,�.�9Ƣ,i��E����@�q����+l��Ύ�8'���w�?*%ɢY �&�c�܁�΂�ط������նθa�巓��LZW-��G=����4�&�v)>:��Š��t���~/ɒ-�I
HRȅ����f���՚�!��� =�~M��24���d3D,�U�������| H�[v\i�2�՞����ѧ��h�Zm{Ě:��p��o+q������Y���Ի$k��פ|����$���1ZC��͌_L�:�KȲ�Dv{3��73�Y�fzCeYD�y�r�ӅL`�4���Yhug��~l���!}Fq�B�`cM��GP?�Ot8����o2�������4(�[���PQ��20�� '�`,���Zg+�0N�ԣ8�pRr��@�\>�vEH9�����-s'	7:�_�L\}�td}9i�n4�B2�y�؂?Y��!��VX.7��|k�w���}`�ǅ�{�{����ͮ��1���m��Y�E#L:�
�@�xs�9��������yh�c���u�<5ÇP�ch;q��p^h0�_R�pB'��=6�ϲW1�� ��4c��.7�ș�M����z� >�
[\O��{��]a��'�6��(���z�h�>�x��v�;o�&u>B|��d�-�?}��-Ξ�`l٭��\|���O�b��t@�Ȱ��|p�6�(�V�z�Pf�� ��:�E��=">�@��v�u�$�nq�4(����5������k`48��AN�!�k��VSJ_iSU�V2��R�ZT��)�#���#(
��M��j2&�7�Eb�s�Dol.[���}��E�=sQ����RT�4O�Eh��:a/�-Y�{���e������k1��	���p���v��3�]�����
��}���b�#mb�3vDp6 i�l��ѭ:d-�!��{�g���F�#q���ƸWcZK{o���bh�����r_��� D��. ����%SX��Y��'�p��*Κ5�K�6�k{k�!I��^���V7D�ok���V}��������ӻ�jEh=(�;Ǖ�O��*�ݧ�] �V�Ǻq�����:���5GUa�ײ��������.-59������S�4�
��S.	�~�W8��]g3����X�΄���̦.ރ/:��/���r)�r>$��5qݔ
.nU\�ݼ1�t�JfC���W�S�K7�t��@u7V��jF9]�*��T����;�(:]�J�R^�h���u�ܜ��V���an�(�$:�"wЙ������يW7�]כ�ͷ�%��w���6�饔��j߮{//+�۷��&Ei���йU�{�;�FM_t T����o��W�^�sUsS9,�����"�SN�6��;Uv�-�9�6��:$��D͙��uپwF���__?�����ϕUUUUUUX�k�[���f}a�\���r-q�v|'=mV�s�	��5:�]��ںۭ�n�<��mM���=��sX/���3m�6V�f�	��@u���m3q®sE.{s,G]���d�x�������\{]��ή��	�����a�ٻb�0���T�+x��Ϋz������{e<�ў DͶ�n��n;,�����>�랹���ϰiϷ<;q���' �յ�pk�Շ�[�_Q���t��9n�`u����۶�n9����;�j�<F��=9ر��f�Q��n�(W<���nA�d�0�����tg���cg������ml���7l�Ψ��r���t�A�N�9Ύ�uw�ώxc��[v{b��s� �Q�$1��$g;��l���h����D]7�¹��nN�7��v�&+<��8��=�6�./���ՠ-н-M����b7�۷vCB�ph�-���=���k7M����2�Wj�n�%�5��q�"�����%�P�/>H,cZ{��v���q۞�.��ʝ�h���콅�����{y�$݇�>m��Ż�ڝ5�+����n컄����	nf�-sv�G��E��a�r�.IG�J��������ln{gb���H�qn��k�_��椆f��o[�5�;)��+m��a��n�X����������ƸK��누8���u�.�K�����I��}�?�>0��]��ý�.Ə8��p��q8��JH1���c�L?!��We���y�z�wL��BZ`�>6����>4 �k^�cM{���V���!�a@�]�m�x?>��Gի�,���L_ӄF	�[�q�	F�pe�E�(;[�`gd,6�m�$܉�w�&(�s��,$n�O���*�e棞%��l��W��Hpc|�1���R�b(ߋ��}�.f�����7o �o��g�Yi���;mA(�6߾�K�)����5�EV��{_F�j�-A��>^����Ĉ��bW�����.1}���Z׾ܴ̍�"���Gv3�&�Á֢m�Z�i_z�t���gjJ;T���6��N!�/�yz
>1��m��0�Y��a���. �k_c�0Lm��a}�*�J���P�H�o�+�g�� ^�D���gܐ�Bm���V_�_��(�U4HCn��8~���?>ܹW��\�ۤ:�0Z6��Ws��ۭw����Zp�w��a�>�����ݠKx�sI�A$��۾�*chV�{��>�g-���N���l4�cش�m-��u�	Er\�<[M�j�#`P��-�9�A$�֑B�ꃼ�z���N;$���3�ɾ�ѷ��bۋ<T[ʶ���h��%$ �6	��:������F@x�K?~D� ���m�3�v�5���
s=�x��3m�"�{�_u�ǌ���F!��Ʊ��_q���-����eǮ�a-=>�贍�F'Zm��Z����V|����\��F�mw_�͵�ܳ:��X3mƃ�'ޚZ��!6���Gz�������b�t�g�!�J�Ϧs�Zpֈ7Ò�b�g��{� M��_�3\�L,M'�8 �m\Pn_����a~���jz���^n�;9l ����v,�^ϴx��"���\z(�`���F�y����-���S�$�<Y#�j��%V��K=֤z����y�_5�y!��;�n!���-El�p�.:Q�N��.��ĹnId���4�>4�s�t ��<�]ׅ�C#�ȰP��$�ڰ6D��Ƙ��r]�p��{�ɯ�D��LV� 
�\4G6��FЌ��>\Q8�yke��,�]���[���=��o�A��n1��4�!	a�k)ck6@1{�.	��M�,h��Y�0o�%A�x��6U!��M}�1gသo��T��5���E  ��cL�f6S>��i��qU���z�:��Y�v��h��7��jꙡ�
�M��=5�-�\�|oc$є�}����B�]Ư�۫F�"_:`���	��]z�,��Pam4	ޯ�y;d�a�ξbۇ��3�vt32Xh�9m�6���Nʱ���l�����<�z�:Xjk�;�84p`������*}�>[��L`�w��v'7PPf��w���c� -p�g�˾3/�^�}�}x���@6�㬶�21ڑi!���J˵�B��'�������c��5uG��Q��30Ё&ڮN�m�ﳎ��r.��%�^� ��#�G�9�eې�8��1���s���p�, Z�mu���b����-��w��>�5k�]���]@�h�d{��؀��Em�y�x��;��W��zkق��#�ۢ�5^ڱ�����>�i����v.G��)��'�ӝ_����H�W�8b�bÑ�5�߷���{q���� m�b��#^�,O]g:��k���'r({Rgq0B�&��epXǫo�>Wd8�|@�������.gXy��Ft�KS�a��z٭���/�g���Zs��Rb��Qh��*���'%�?/C��{k�QQ6%r��E}�-Cy�|k�N֋�(d��Z6��Q�������tF�C���؍V�2D����%��3�ӛ���b�΍h{0��-�wA2�cb(�q����WW��Lf�ѿ6x��u�X�謋�A��y�tY�4=���+c7-����.�D.n��Mղ��h�!�Q�0��a����"�#���rE���pR� �L#a���g�y}]��@.2L�@ |j W�h�"�v&�@��O_�}b���@>+M���\�'f�G��C~xP�1���N��O�{��|/��� ����CW�+3���FY�{��F���<���A��5��o�oZ�_M����������d}�W����hPhs�Ú��{5�`�6�\���˟}�޴�7ε��<�0k>���E��
�Y�*0���!8g.�nOZ,`Ӈ3�-��ȁ[P`@����)h�ӂ�rK�;zm���ĝT��H�,�CAl����3Dw�cj�H�6�R`�A��C���7<g��]���R4�1B��C���?9!	��5ac����B)S���䅢C7)��6I9X��{y��4�V�	�{�.��J��j���^�*r�L�<����*��ܛ2U��\�v�m��*y�K�ƑH;	q]����LA"Օn$3�׽��zR8���ݪP�BsT���3�W������f��0Y3��q����۬��%Q��b��vw�"��=\�7��j�vz��{����n9>��GBH�dck�L��2@����H��!Y��"�q �~�-��'B�_~�ߵΎ, Sx�� ��+,d8|�m���Cl8���ڸ��$[��11`�
ﵨ��q��o�G������,\��+���n�K�bN�Aw�w���{7����������C��L��Pa�� ΢cL(;��˻�����5��nk��w,�E�_,��A�)�e�jvJ���GţLj[�9�p�u�e�8�Ԉ#Rx�^�Pn�,�D�3�t�<����h���Xc`6+�-�|M�#���W"�L}$�V+�L��;�6Maߵ���2�@���x���]��'PZoP.�k �y�Ʀf[�X�ZdB ��o��2�-iA��-�����blnF4c�O�=�g9٧5�[&�R��e�������oO��n�9�֭J�n�[k��X��$��ᦩ�QFR(o9.(ޡ͠F������"`-�B@��u�i��-s� !��Ȥ;þ�������ϸ׀��"��0J���v�rƞ�o֋E�Cx�d�j�&��,`|�{�fQ>��{��󫆇A��"_�ke䆻]4�|'�%A����i�8.�a�[��`��
��@�"m��s[El�2�;�X�:���E�N��hl,�?n��V�j��ƾ�>�aR6��|2qɭǅ�E���v��E�P� &�w��}���ߓiк� ��F�b}눱薙�Y�b��@Q�тh�a��{���%�F'ִtЧ~���}�pZ�˸�1�K�Op��"��������R�0z�~&6b�w'-�x���۲���� &P�����.�ڛ G�j�!p��t~oF4��c�Tw�)Z�.�Z|�?��յŦ��sB�.�tP��k���c=�A��h5�U-�!�k���
?x��P�d1�sX�L��\ɑ��۵��v�zQ8��(���;`�~~>B�+k����������q�1����u�#�����F� /=���E՝�_L[�kR6��(����vV�m���1yw^u]��n�q�i+8�Br��I��KJ��y��B!�v�Ac�(��v����e�tA�	���b4|��6����t]��{�ܝ��(��^��P]��X *4Ռ�$5��L�닆��8�,nƘ�:�/D��g�@ë�o��[�.gi��ӵKu�ѥ{�a�~\��U2�7R���k���\d�`�%�f6����K����r����)�ݿ��мs�X �����I��6���v�G��<Mmp�'��Z.9���!|� �6�6���J�'��E���x�|�F�]4���'L��z=~k����Y�m"5#ѳ�0�_vx[�j��0���>)�g������b��%|s~v�n���!; �B�m�O�_{��=�,�h��Am���j�]�w��F	��9m�q� -w���x�M�K�Y���z-��z�,����D}_�����DYM��;ܕ�� �9y��֡��/{"ዮ��y���F6�@�}�z��
��a��n�(}�[��c��'F�ȹ�S[]_AX�,��8�jJz�φ�z�8r4�Nf6�d��±_�(lr�f�A�w>�?n>b������k��I�9��0���[��6���/G�#�{�r� �6���e��Ώ7>�Q��6�K�	�$� Dww6f���a�gUݞ�ϷYPVBX��(q������Gu����v�E�q:ର4y���p@ߴ�}����DNE���N���z�!�� ���d@���08�;�V Xڛ�w�#�,>����T�7��:�V���a{C��-vzH��~c���d���mѤ��$���~����j���KD�9��ᦄ������㮜:<|�6 �~�Zt~̻dȢ���m�_�<t�s�`P�P�D�������>-6<�&�y�#}=}n����Kb�%Z-Y`h���E�7e�Xt���Vxg]�@�)�����V�Ѷ6�� �'�G������Z�F7B$s��{��<��V�l-���}�D�@  z\N;@�w����]���A-�:�0-�/���h7����\P��y���5�m�4�:�Y�B�o 4y���6w�l;L@��O{]c ��h9�y�����@><L|ۋ�5��|jK�,1F�Ek�z+�~Wz0laq�o��ua�$�M��j�DA��x��֏�~�e	��5	KL��4�`�Hh|��%`aJb��O/3/Y�q� <S�a:<�#�=���n�K=�y�H���`��}땪e2j6�w���@�Ol��Dա=��X46�䂹)DQ��"��x�k<ӿe��F�DO�Loq�g$q����g��~'�u���m����.�v�YHq7	�x_����5ۚ��y-}>҂��������Y�u�bF����� ����_�_-�Q�;K�Ÿ�]OK���Ͱw[�ޝ���k�;mǳ�v�8:舼Wk����q���
=n��r�b���,�׍z��p��X��g</if��l^/X��Xա���s�a����f:n.��w��9��mܱ��N�Dfy�۳�tܓ�����'���w�oZ��p��8XcJ�"�bۮDn�;�x\V	�0:R���Lp@�Q�ղ&�x�<��/k�qo�� y�LZ:>ߛ{����j�H���L�Zڲ�5f0\m�(�'Ƞ`�x]�(!��0t�;Ÿ����
��_Г�ǌ"^�8N�ll�!	���3�i������`+cN2�G�r+2gc�`�a[�sN��1�Zat_b$pe��>v��72g��s�a
m�����,2�X_\���7������=S��d�>���G8�Zt�x��"�:h��sbNI�mY��V��A%$i}sB��ή�>�lSքmi�!,��W>V��xkN䉍q�Q�H�"�`K�;PCl���>$l�9�>G��w�ְ@6O���1}�"��܊Yd�/r-�-�E`cLE��o="
33o������=��O^u�"�v��/g[���Ƿ���|�6����ȣo���5'�^�6�rɞ�P�?�H=��[�|�4�1�da6H��.�W_��#����=J|~ ��D��دuvh�\x1A���$X��_�$�������lBέK�/��?q���@�u�k��ef�W��S����R��Y)�>�%�ء:}Dm= &v�K���� 
��Aئ}��6-2x�m�$�;�M�m"I�������X�ʠ��������bҶ;,���=����>i�|�ֺam0%�dA�����ɗ����
����m���D���vѴ#��K;w�M`�#����	j��T���쿙�1���l�G �Lo���f_��(,�2@��{}n��Ƞ�Ծ���z\�]��[bq����8}y������]+֙$��R���M�vӔ�+���^�C3ы�u��ޕ5�;pk�֎�Fޒ� �A�[��˲�)ޜ�1�L@������[����e��n)�m�s�����ly#;�Y���:!J�.cP<|�s%�bjr+�`��s�o��_c$N�6C�n��<�>y����Rf?B���|X�8�MP��N8�"F�.]�Q�*��+���'��V�w�kڱ���&������֮5f�fLr��Mp�3��d60)��Jay����u�K?��q�p�F�}9޲'j[�-�����8�����ܼt�r�'�3���-�fٱiG�|��k��+�l�If�r�aʽ�{v��Ԍ�ܻ���f�8�.{�[-�SV�]:�Q��M�沩�_Vo'\E���o'^}ݗ5�.��Xs_uwl�����mA�	8#]j��^�곐,�_F��I2�`��RtV��c\dpdq�����yB�g/��͢�����3����on�=,غ{T��5�!�P�!Js&9����gZ�N%t�)k��SZ��i��D5����0S���C��L��;�._)6.k��n�����ыS��xo%sy4mmx8�c����9tK��NN�U��$�5����(�gwz��k�ų���.��z����5�%���3�r�u5a�]܋��^�k��f�vd����S�7����D�г��=sG>���J�F:rw2y=�|�V1j��l`ǝ�sd��w>�u�j��y.�
룼��t�+H���n���<j�����~��Wn	}�@��/�x7�;ӧ�*=0Y�=����� (׺��{��]�>�p5��%�|l��s^�Mq�\\��5��k�Yk�ϵ��¸i�ň�t�b;=�����"s��ޒ��	���G>ݏx���,h��n+H@���hm��P�131��'��~��k���v$aP�ao���o��E��ӌ�Y0gg	h1�����$��L������)����2�dA�����i���!x�5r�P[���
R�������1�}�^)�婖��A�,M�\��C5��7�繎<l�l��B,���䘏1��3�p���=�N�U��vwZ�[�'�H�ڱ��)G�|�;��"���[��Ŗ�>9���8;��Ԍ=mTG����=ǠN!Jv�������Z�%�$u�E�k(rڂ�ۖ��_o�}���K��3��Z��]��r�&�Ť�_�׭��2D"��%�`���6�J�s_W�rrD!��^���n��&�(�)�w�*S��
C������ ^�����)���pε������Lt���FX���;~o][w0x/s}�/]�8^[R����+h���t�JI@���_�h��N}o��,@�]���=6G�ق (/��c;�Gu�ӠG��R7��cW�y��� �X
�������I4C+��W�0���a��DB��t]�m���ω�!Nr�#��nGY.n�n�a��n�q�:˻��>`��-i�����4�;A.AN5�v#Z�i����X�\�j`(����}!Z<�B濛�G�|Z�@`�m����C=���۷�m���E _d���On˫P�'z�G�8j��!:�24!>+�]؋����ϛ�����+_+������i��o;)rF��jѕ��w�.��B��l_dS�:p��� mNZ����7�4}][�������l��:\~|�`�1L�>!_SVUƯ=�glM;�dY�o&�Y^��><P������ �6 A����>X���x��Y|��� E�g'9CDn���sz�	� ���:�k�q<8|�ywS��{�R뀣IP���M�/��[~�h����&�Ř�k�;^o�����Ϝ]�����L�,�BG��6�@�w�E^�<��;f�6�}v�|�<�WJs�;�9x[�4���d1����I@B�f�OW;��^ݳ�ɘ��)�]�0�n���eE����/�[��:�k�|�|��v�7c�!�қ�W�]J���g���ո��)(��v�G<&�n�p���ڧ��O6�k�ܞh�mح��x��\L���H�3�����G�GΝ��3�u� 3f�b|ub��� �<J�3K�k���k���Z�& �r;��i��^^��d/S�d�4~}��#j�qz�0�e$9�)	��m�0��y*os>ƴ\��Z�u��x�kX��=|ӷ���^vٻ���ӫo�C7!)Ig�b�kt6�.$�q1�ܔJ݋p��x��9�i8;B�&��O��f���V\��"�Y�>!B�����N�#L�.D3�!ik�\�x�����YlA�/3�b�>)˲�;i�(����b�Y���"}&~d��������o}j7���i��-}Ư���p���V2o���$W��΋�Yȶ��_��h��mf<�w�<�����5��F�� #����4�\)>5=���x�� ��^�B ��E~����ϯA�$s�ݺM��dݶ�f��w���������¸W��0�dN�hш̇�5�tG�e���H��p�SG�r��]4��`�����m�mGf!s�����d��e�[&-3͐v�e�~Ư���#��iN*�k�s����Ȇm7vpO)������*���v�<.�b���Pk�:�=
�f�Y��n�\&\��?�������� Պ>��z����� �2\v9���[�붲��!�Z�š�m�I�ttY���o��=���Zq�L$��ݹG�0�O��3H�^�yÅqj!�4� �z핼���j��h���l���tq�2�*�����=��7�qi��`��J�p�;{)����d��<=l��]s��o����߇w_� ��s�-��־����6j��>��6ch4_X���\�]B$^H�F'�Q��Hm-h�T�[�)�Q���r}sơiF&��*�~z�IK�A����������r^竄	7ۙ�q�[��+�#�qS"�XȮ��G�a�i��z�� Afv��=4Vct��g�ù�E`��_ZX ڏ�ᆿ���e���_\�/�qݯ4��m� ��Ys�q�qlB��s�a�p5XX_c�3$�.?e���+��W���½��y"�#р��n;6sfJ�bF��B� �H��țm�l7�u��M��`����VkN8p�80oC�y7�|�����!�S�o�ܥ�%R���=�`r���ܫ��ҏ�������Yؽ�ƾ�
c`/��c��}�
GX�/[�cv��Ԣ�B||� �j��Ű^��Ӻs>�Ab���Y|��2_�.c�ayp��؋j6�܊�`�2�Bu�]�K�m�0Xtv�Ğ�{  �k�+� ;�іb,��{��8�扈/@r0�hA��}~�{��o�{n������8ȷ�O�D[gE
�ϛQ�E��.o�����W��{�Yp�D��ݴ�-�mZn��ܧ���g����>H�kL*���NA�s�,(��?$=�~ԉā��:�]H��事]�N+��ሯҨ0P
�dO�Km�ŋLx}���^o^E��g~z����$��m��޿����]�i�����]��<�O
<p��&z_�����ȴF�4���|'�f��P�Kݝ��O�\�b$�1K��L��6�A�,�5�{�V�o�PA����Ω�i��fq�z+v����s��`�ŝlL�}o���k#��Ƹ�W�a�;h�Dq֬m�GG��9�����͐�>7Vg�\n�L���~�,a�\,�����<� ������2r����nk�r�򄘖Wtۮ��vi�ͬx�[]���c�[��f���z^7�#;e���A��^��A�����4gg��7R�Q�ۅ�} �ʲ\A����%�g'�yk��>���F�i�7�)���=ƹ���~-Y�u��Et빆[�lB�����ڌ�4\�#�Hy�:M���j�n6�x�m۶ޏ9��L zN�g�2M[��]��9k�F��D
��-gW��w�
��r�Y�PЎ����^4��A���c���9bq��w���sZ/�u FY[�77's�� +��?���IW��1۱X�^�/�U�lG{�VXo��|+��-����Ζ�7d��pL�!}p~@��B��A%�v�;������j���涾0ZG�~���g+����b気�A O��dx٣+��-?��4[��F�=O���,�!r���1e�A
�|Q��\ƸUЏy�d&��O]�����\x�$d#�v�N�\���Ôtu9��V�O�fog,�,c�]7Ӆ�b<1L�P_e�:�r���(��a$}���:��퓺���o,淩��\�3-qܝ��WC��ۊ��W^�}�췐�$A�L����oV[�wD9m�c��˹��H��M���2�%{tr��qep�u���v��k��v�e�/M�ֲ�ۯW��wo�g-ύC8�v۶�_���=�3�ܙ(���a��n����^���Ie�Q˱�Y�����<����V��Hy������;k�ܤ�NZ��,ꝸ#)��uȋ���$����m>�s�x`%���M8�U���1��P�n1����[�����TRZ`n�8K@�_��7�+a�^�ȃ�̖%*�8hIDQ��m�%���*�V$��1���_��4g]ڱ��%�C|��\�eٛ�)�^d�\:>ٽ������LW�%�[ ��Sp��!)��Ds�7��HO>�ɑ�M0��b����\t�Hg�Zx3����`��I���^j�uO*�fi�<,�3�E�P'{y7=��־�YW�y���x�.�G��>G�-w��*r?j�~<����ٶ�κ���Z�zͭ,�0��:]�.�3V��!9�S/��ͨ 9��'�n�o|ǳv�q}�N�]o9����Rk�>܋$戳>�Eك|���$�F��54Ԑ5LXC�\&����,��E ��	�۷q� �O������u�������省U�l+X �ל���"�Ű�uA��2������zY�,���=ss��t ��˄�����\9c[��$%a')ƽ�-��70��^>/fC�uxF��.\�3z&�_�̾�z�J�r!��v�z�O<�N���\2���ꖶ)r�Ai�<O��3)�D%��3�L���Դ2]@��Ce;γ�H��,��90�*�z���$ϔa]v�����.�A
vpVE0s�z��lo�6YY]��0 �Z�p�)]�^뉋�K�/_<�ȸv��ά�����-��a��0�:�c�7�k�8g�9��$7��S�Q���im��!凇��e�8�k&s�^�Z�1Ԏ����=2�ad�Ljr ����U"�8�-*ľA���/l��_vx�%]��8�y���O�}�B������^�U�Fp|�f�C�g��1��'H��Z2fK��-ߝ�����{�O��M�#�ǌ������z�?�����{�S�-c�|�h����X�����6E�>Ww���דu�̜��|r�J Z�Əy�N�����X&�s��A�VA�Ŧ.����,���]���#<����3Y�y}���Ǔq��{:�P�Ab��v��5���n��0kۻ�7�ܚ̓�b���ˊ/=�w%�cU��>�r��Gz����#4[VR� �q�س�cX�c=�_5��8)^S8�g.��]�<M0g�¨��=�\��L+�w.�}�(ϊw"PE��+b|�/O8w�����"1���lڂ@�O[����`酐�#)Ûl\Ļ�uf���AK�I�C�r>�s�t���E�h-�`O��f`9R�	���-��[��?L֢X)�cY����ʷ�rİ+���ƅ=����jۇ�� �jq����	��������-x���F#﵇�����߻4EX�f{�����B ���iwAUμ2\y���5��]���ꚽ�;-\�6�0�V%;�v���k��$�v3ݪ�J�|y���&��w���p��%]YՎ�_��!/3]�[;ϯC௯�+��W\tS��eR��YDg>��w�nór��qW�M��=K���KC�UBG;��_a��r���Y���w֔��7x9_6�0���"�R��a[�g˻��������h�<�07�uÍ�=��s�NW�_;��Lp�^4��g������귴uج��oL؃������ne�y��y�S�Ok	e��3�/O;wL�r�z�_j��v�'9���iTN����|{&b��$^���	�V��5�w7t�ƽ�l��4��s�79�O����l'wzA��H���N�^q�M���}��/ke��#ru��I��q%���2q҄ݝ��&��k;)��ێ��mF8��>RrQ��N��_W9|o�n���w��<2�wt�ޡ�����I$�I$�I$�I�;�m��N�,)e�ܮ�Fzn����q���ݰ�f�A�d����Z�<��q2�#�|��K���0�p�F�p]T#����O!�6��;�r��4�[U��y��1�i��䳯%�j���0��le:ݹBwgm�����K�{i천<����ð;a��b]8���l�4�n�nK�n��t��c�V�U��-����ܶ�\��9�v�T�Z1k6�\�ݺn��:��ݶ]ȩѷE��<4n�}����7=j�<uS�v:�=��\]�����Mt�ڻ^�t�vp�8��&����m�:�r==�j�B+��mٮv˭�]�氙d &�iL.���:(��U� -�xURl�;P�0qqs�c�5=ln6��9�=�m�L2���Zta�[���x݊��ɶ{vx(�m��`{R���BN
5��ɸ��F��v�ۍ!�r��� 3��:�.ݩ_l�AtG�m8�s׷���x��u����j� PݓlD6�!��Ӷ�iw>%	r���!٧q��v�:y���x607W$N�e�?>z�_{�>���Ƌ��.luՍn$g�/j����j��]�{n��/�r].�w#�D��TyW;�������{�<�����	��c���aէ��ˮ��Vx:�c���6��U9 ��w�	��cF���ۿ�O��|����p���$������\��vZw�����Q�
�۳B��<�o��޾�x�����f��M� ��(�h3��yz�������%gf�N�_C��l"\@��WK �̅a�&��&��l��v��;1BӅľ���΂�h�x�2V|J0���WZ|��K�8׀���o�^m�Nz⅍x/`JgB�xy�~�7ڼIy ��N�"�Nh�]g�v=|Um&��;x:0�	��,�@�I�K�*_'���ue���	�j���Ǎѕ;Ub��!u�]����"Pv�Ӆ��r
ǵ�{)��<�f�1�4J���1e��Y�~�\hѾ9ia�l�Uz"3fl��{�9;A�ǰL�6�<�F��	yʅQ�in �����撚D�4�{���u�s��S
�4`��tk`�� ўR�]�����Ó\�ڰzAN{�Gr'؜�ik�>��A{d�#���TQ���%�,;�N�جb�k/��O l���B�|���w-���v�<GF���t��k���W�P>%��9̾� l
��vE�\�����Q�I��;���00�9	��}�a�]#��0�X�}�]�b임d0��d~�c�犙
?fg}�r��|�J%	�?(��DS57g78y��;�p��_X�E⇔u���D�ӺT�P���e��k�[�}�+�]��DX�9)�d��Me�wugt�K{b�Ʃamw$��3w���Ӗnܠ'���c�#�,���e�=J5;I5�T��/��u��[ܖ�Xu��s���ݚ$���Hp��:��N)�b�ASdś�	�L�i<�I�lZO�̓��n��][0����Ϲ�Vmq�kF(Yc�A`�F�O�#8��.�"�Y�pba*���y�1gO���V]^h��C�G�c=������~�����Mc�3/�؞�GZ�.-�]]q���~�|�n�5���e87�6ҳoY�P���l	M��ĪVM�c��>�
1������Ҧ���E�nƻ`�!v�Q�ؔ�|�Ή�i	]�_�OM|-�����W�����ʲ-�=xS�����M���v\֏��!<S#z�4TI-?=WG���=�x��I�{�4%���`��J�w���Qc��Ӟgnࠥ-��v�;�7'�^.ؕN� Kݢ��	h������@&|�E	� =q&����v7���Iu[%
'`�ox��x��Q���g;:�p�%V�H���$�m�ٳn�ÈUkM�|�8�-A�'-T���;���ƌ��V���`z�I>-��Y|ɻ�b[��93)?�3=o�����̔l��^�* Ά#��C��N�J�ϹJ�H܌�b�4ov��8Z#3[}���P�9p�2W|t�#�"続i����A���6kH�
�3EYv����;�X��xXf3�4��[�'Q�È�����99Ś��N"0�W�� @�)��wL�r��l��p6	?75N���7*�'@�Z܌Ӟ�I�k����z�:��r��۝�N�VV�����h�K�Vuo@�)r<��9w�g�v8�<s�b��Ha1ü��=Gq�/k�@tz��s��2c��&j�^NS����<v;g�g/f.ܨ5���N��&�y�v�A�`.fփ�ѕ����]q�O�u4U]s�s�)�k��&'�ݾ'0H�xZH��Orc=K��G�:��zV}	8r�v֮�w���ϼ������������)��>�rPz��-����E�//jzL����Ƕ������|;�M*�g���y�ƛ��㌵~ME����ֳ 2���Y�8��vA���7��R�����Y��2�a�����Pń{AΜY�V�н�"ՔY#� ��C�:�'ș�4}ඇ^4*}�	�Ҋ�6}�r4�$�"l��Du��*�*M��|d��M�uȕ�V�u^ 7�,�,2�O�0�3���ཱ_������G9ˇV>ukzB �3v��G�w�q�JG�5z�HYϗ��ے�Zs>���LJ���b���Q���r�ɷ�Z˔5N�CI{����N>k�x���G�*h���p���t�7A1 _�Eۖ���c���.����<��@t�%,W�����i�e�|I��lL�a��0kȄ8�gU1ބ�]�&A��p���츳�c��엠��gM�a�v+�����Ur��[�kDE�G�h͜z10�X�"�C\ힻu�A�lq�a�� RF�e��]9�1HIo.bG�f�-��Ȱsh��fôl���d�J��l�%�AܘH�q�_�̩= ����[�����,�,לZP���}70֊�k9ϴ7�/��ڠI�����M|�e7B����W��w=c�N�yb�0�Ӛ�1�������Z9s��Y�j��{!ݛ)� ���4tK�ܴ�7'N�D��ƒI�h�f����f�V��Ϝk�+1��O���/D�6��izN����ch`v�Dۏs�3�7�JX�æ��ۥ f|�z�`���3�]ݺ9G�?f�vCc�8��;d��nzr\\�}/ɏ�=��!ѹ
�}�^�k���G�2�tzL���Gc�DVx�䙐�4J��d_I�� N\8=����xil6-n�yn�$/�6�*n�Lc��1�p�ĳ��4�ٻ;Mn�epM'Z�xJ�+�2o|�.g
d ����{I�6le�}ݩ_C-�����U��T�������C�jލ�t�e<;�]�Y[��n���/L9��^=6Yע�Zý/)�L'g�r?��q	�9jkG���v��h����09��Cn[ͮԝ��˛cmYV��Û���-���`��PGn0�c�6T� �-�ߣe��i�0e��HV)*2��j�R0�m6��@�~��Q	0p�)�rf�������c��X����	��y�c0��T���#N9&S�+~���S��,M�Fy���O���w�8�;��9�;b��3͋[i���DK�az^Vq��˽�!�8�a35����2��V���׸"�✃��Ԑ�:�����N.�ofj{�a���y!�%`�R:���_�x�>��01n�;�gk��]�ܑ`���+���d����I�͗��v�&��q��:6뱐���;�m�z��y4i�T#��K��g�pv3��W��n�e��!�N���6ּ]W��M���`��\F�q�;٩r&��i��8���Yy$�1v�=s�W�m�Ş{2ٸ��p��n`�A.T��˃z#�&!�K��{�g�f�3��Ӱ����fN�-����
�n�� ���u�����`S��ܨG	 �nnns�_L���q&T]��d��]�%� ��L�����"�ٻ6d�ѓн�*���2Zl��tcy��n[��G��&�*�R�Z�3T#短��*7�ֳ��X�O4�gp"�3��.Ք�,\7w���$�|4�X�ni�L&��ۛr$�Rx97e�S�7<l��PH�������/�vz�wJX�P�]��$BR���H���\�v�/J_~��M��,pOtW�/P���m�j�'��*�=����D�������I��S�aⷧf%��ڴ���{y���9/f���x>�=
3����n��������K�*-�Vô��{�hI��e����^���(����G0��m����;�ST �u;��l!�>�p�2����_i��uٳ~y�Qķ8H}���C���ut�g3�q9$r�P�QoI��-�s�;Qpv�����!���%"�m�8wn�<;)�!���Yfx둶^��]ˆ�z�<�id�:Y��w�%��cB�i;Έ�gv�MV,���U/��׻g��,傐����L�6��1����M�j�q�v�X��E&VnA��@߾�/�~L��||Rѡw7+{B��x����6C��8����h�����״��6���N�:�~ݎ�[<۔Gםb�-�v���h���Y�����J��I�5�*h}W1�K.��~��o9�ή�5K��Ά�d�Y�E�s�L�E�Qbqq��m���3N�������mW���f����C��Q��'71���ԍ�>-�S�2ള\F�#g�ݺ��d��nu��ˌ��#�d"�>����:f�|�<�\�C�����AM̒��#R̼}Y�<[x�['���6�N&���]�bXΊ�W2{2���
c�������6������ԫ�m�=|j��7qc�j�^��M=� B�/L���)�Ծ�;�;%	9q�u�5�j^*W*�#����X6��G߶�,���2�\1(��:��7�<i-`I�O*Š�ܽ�
��t�>��`�l�_�\��u%�e��g90��8<O� H���K4�28��Vj����>�ѫ�WS��z���l�=��Ph9'<�NL�!!�.�aؓ�ѭ�Z}�����6��T�|aa]����H0��!�����š�>���{� �H�8���Dؒ��[b˅WH��R��o-�e=BpI��J��#�3t��)ͮ�/�fL+�*�p��Ii�y�K���J�ˣ|��]�>w3��0%�W
���HN�z K<��-�~���.�i�{1{�}f5V�v�m���y�v�U�՜�烽v#J�
yod�O	+��"X/���[d��rz�w�)z���^w��0gwb{]��m���od^�;��	�;O��D�ڞ��N^�3�ɄI��;b��WIiq��,� �Ϊ�:�u�Z-����7l[�-��RI0N����ӂ�\!���f��U�&��FX�{,�n����d�r��`��K�`�Ա�}�y�;09[���4�����U�7�"�N2�ㇷ�4��T&��O/m��ׯK�j˷4L���Ê��u	���Of��Q0���7L��0CA�O1O��G�i8��nN>R�Lf-\��E��Ja#tf0���|%ɦL^����Ի�k��hx�\��E���y!�W�Ѵ�84�E�4p���n����ɻ[�����G_Y�ի��.�8f8�FM�9�AV����v��x���\żKnS�=J��Eݹ�qnm�;X9��'b�H�uP�m���\nٞ�]۹�7`���"�3�� �>D���ܟe��֫�Vxfǁu0Dt! ���qCaU(`GR�}���aHF�(�o�+��h��y�F�ʛk;'�vD6��ˑ,�u���������w�Ĵ��v��#R�%3����>/&x>:%�8��Ϙ�s�%��cvϖ��6��I�o:5I>� �UmV�<S��x��#6��:�j!�\�QX$WxKlw�
��IF<Q��zl�R�7p=4���S�cI�oC��n��g���)r���4�?K�=�z*l�"���ɯ;��ua�?W�X3H�O�� !��b~׮p���s�R��bQY��vi}������4%W��D_'���f�8��c[O�୥y	$W�2��V��̱Fj��k��\�!7&V2g(�z�̣ ��OQc&N�\F��;�:�ν͔H�d8�eqk!-�Ԩo�ZCs��^�a�q:l�y���j�,uVW13�k���h���Wņ��6wW>ݾqn>'���`�ShR����O�/Ϯ��޾�}~~�)]���un��O-�t�,�Ύ��M���!QJ��n��]:%�ٸiu1���C|��1���\8GK��8M��0�59[�к[nj����͙��^��ǆ-�C9��|��+K�DuUKdP� �M���g�"�E#��w&��� G�aT{�9��gm��j�c�n𮲻]��uj��~�!���Y4آ|�*!�]ǙI�	E������ksM�ݼڝԧ�/�vg��$f=֓��l=���\>�������a�{'%`������Aΐ��潑�r����P���[������??c}=�*a�TK��Ҝ�;��9�P�$OϿ���{��vZ����&x������46&y�6���ϳ�	3��#EK��C�^���c�� C��n�x�6[g�Ũѧ`ѿn7��ɩ��܃{�v�r4�41�
������gk�ԗ��l��G�x&Fo! g����:�����z�^�<���?&�}�.�i���ݾ�7�j�*�V���W��R���9'��|7�e�s(rS.�P�ڦ@�t���	#�&��5b�f�}�����t�7����˶]��:����c�������]�G?���nك��9�+��Kea)6q��L��i���rN�.�J��6�-��9��_�cY�qm��C�Q-h���q�I�ސ@س|}`�]q|�&��E�����-�ü��� 
�-X��d��
6=��b{��uqE�>$���G*��sIc!���Yv��m�����u^���I���$��z��xrœ��QIv"	Pe��4��~��ymD'4�I�}�*^��q�$)����}�:Qff�P�3��5{L�O�5U띖S�"cf\�J�����oϻ�������)ޫ��xV�q�9�!�[�N�1��5���4�s�sZM�oq�:��ü�i�#��:f-�qu �i��۷n��u�"7<����u%�|v�m��м&4��e��SN�\��&�]sd���ݩ�:���.1]\������xO�C��Ρ��ѻ��}��O^Աy����3���Q.y��hg<w^2����S1����_k�-g=�b�e��N�niĬ��,Y���{B��t+�[PUd����4��
]�{壼;ӟ���tA����$dL����!d�↑�E#�7�WY(�*��N��D�=H��]3m�zZ�}ՠ��Y>�6��s�6����M]�M2�,�X(��Ƌdt܁� �N~ab6�#&;��m����U��� �wb��ʺ���ˏM2�	�#�֍ڦ��,����ܽ=[˞&b.R̜6��ɬ;:�±����'s^!�-�Iʹ�F*�Z$��bW�<H����2Mz�A)� �|{SՓ QcibqC�j�r���G���r�I7YB7�x#�@�=e{qa��c;0��V��Z-�6�c����/L�F��w>
���j١I�8
��yD�Ef��l��qWj���:	�/�z�h��r��E�Da��)!�7lrY,�����;�l\,a(!2#�A3��+hԣ&�ô�.����<��J�5ֲ��p��!#>f�1àW�"k��u�`��)�Ӧ�% ���/0h�&�[֝�/�򙩲��y��\��P�(�z���yU�?R%������y-;�,�v�Bo�=����U+y���+*���c�
�v�<bd;�>s�Z�<X�cVS��D��;�ج˪z��p�F�۶�;:�r&�E���7��3"���G�=U�^��w����������V�7�q�[5,�9��M3�d2ͣ!�"")�F�����vH���V���:�su�F�=�Gzإ��=QZc4K������n�[i�uڥY!2���u�,k*�Oa�8�l��З�+9�E�+��s��ٝ곍c� ����Xce,'H��ݵӄ��v�R��¤�%Aw�=m�C9k�˷���d��՝��u�Y6C)�^��cF��Û���j�ú=%4��������V�t���A�8���s�%�g�hz��^N��.����Z�[�)Ƣ%��Y 
\h۵�����h+�￭�w��x���S��)�w7�����:��Pq�+�D�P���8�8��r�8��5)tF�9Ԟ�鯬�;+	��ù�QB8�k�G�6DC`��/5��\�:�/���ä�"�w8Ƌ��3�Tz��	I{�B��v�Ba�S[�9�;V�n�ݛ� �aްBR&��(Q|�>;�e�gq��L͇EY�*�ޥ�e��o�Y�;F�_����wg�%�Q����q�U@���h����޵ӥvP�w^L��N��I'���K�ao&��1]����&6/��C���|������W�2�m�K�g�t�U��:����I;2֎=�T@N�T��q�{O]�ǋ�ɨ^��μ�j���a�݉o)y�]��r%w�R��������ّ��'�P�6=��ͱ������zk^J�/�5û�
���k6�uɿWx�_7r��j))te�ǄV�>�#����P!U��k�z$g�Y;J?n�y��+ ֮V��k7�U�Y�����%Vi7�:5�≾Xj=Y1m��/,����v].o��Sw�^
�Z���.�vViX+�7n�����M���{M�.nF.$&�M`���0{���8�W�������-G�F���ߟ��;�������ꪪ������X��;G[�����x��r�|hb�͗q�eu����3Sr&ݗ]��kY�"�&�c��9w�C.�x�Łx���v^;\�=m�i��;rŒ�L��G��zv&��p>S��,]I��ɭ= i7n�<��d�m{u{E��g3�m$�<vC���N*-[��j��#s�n���n��cIu���۷I�p����k���<J�bmN�-�&:ֺNK��r�ҏ�9�rt�㌞fWkM�;��y����55�-���q]=��n.c��xѭر���{n����{O;��'Mv�ٮ	�r/���|nޚv���F�\Q;*�T��z� ��������t�O/!˫p\4�W2�!u��pc���;�1'fv璖-�G�V3���ɼݟd��l�l$�ݭ�g�
'�U+n�0{�8	6s�"q�pt3ssF.�C��y,{`����Z4�v<f��#�u��;u�l.�mgxG�En��t:��!�е��!힫sv�6��]n9���N:��mg\�#Fm�I�@��b�I�c�؃�S�;&�w�����������.=�qG#Ɍ���q;n�s��ʚ=;�Սn3k{!�g�sv�g���� ��J����'=��7�`���]�v� ��v��n�ۛ6��ۋ�
��։W�:4;�7g��o|�Q�دWn�N��g������r�X����b�������z���Ze��{�"K�q}�r��0k`���H<�����P�������E��1�A����4�t�H�&1C>w�SX��J/�S]��*Ѫ�xQ����`]�ɉ�'�I#����ns����g���u�1���h�4Q����wda"�B�C��Jgcu��u�1˸���|׌�NxT0#��O����~��sl��1P�n0�!aV�b�q�<��o��B,��3�#�6\�\�
Qs�/�D Nտ.'ŋumFN��=�ه�]8D)mտp�ɞ(]����蒻��R�0��̳���I<Uaw2	f\7j�F%2�E�3jy���)	b˳����仺�p.|7m=�!a,'���7�7D���.5������bp���^��T�z$�Ä�1"rj^�8͆�&�y��ΜyӇ�t|����+~o��l�j�SW��*v�g�MJr�X�$$V�u52���#���9�|;��N�g
ײL�Vޕ����4^�(�!����͟4�r��!έ�qEs�v��u���V�a��-`�� ���c��G=9�4��jþ��kb46���{ꨐ��z`�<Y)�F�F(<@(�/ci2e�Ƭ�k�M�s�v�+�џk��n�<Ӈ�6~�Gs�0�����lG�]Q첦��n�s�,�~���c!�r�~��^��������3��i�/ �����(��ښ�9������o����y�y&>�����k���6�����N$НuO�"�{�=�W/�����<N����B3m�F�z��QW��xH=O#7�ɣ�'���h���-��BI�{���ֲ�<�u���R�ڤ@��X\��ĳ!�Y�-��m��K]�Qq���V3�1�lۖ�d��;�)����ޒ�\�"�/��K��!�.;9�����<Y%��hɚ���|_|,'�A�p�
Z�no\�sں�j��z�-�+<��v�3?B����sp��\�z�ݷ���(a9�*`A1��{�Ć��j��ث̱ef��.�H�z�q켯���Œ�3J������L�B1{��48kݐ.tD�p�iq��1��3�������lg�K>��D�����a��s�Q��+i�n�4W�$0�� kky	���d���s�me����;w�f�̘����{`��S���pv\]y��yA���)�:�ySN�H��)���7n�:����ۜv@۔N���sK��|q��$a����m۲p��ֶћn/1i=��D׃:�F���z�d�[Y�\��әk�r�[^�mϤ���\ɷV;k�mp'B��׎��x�`.#U$�g[(�b$e�L3g�z�\ճr����>� Y7����#A`��R��e�eÏ^Px�_gp�=_�H69�C�������q�TEۮ��;��+*h�ډ7��p�Q�	�˴��½��^�r���_l҄~��Y8/�o�����be��F��r%�����䎋ź�+u�jI`F�gigk��ns\��ۼ��;k��j&+��!!�uq�L]u�{D�9̙�P�b�&5�(��Ts������e7H�����!B�&�,�p�C���V��--�ۅ��Gb�f4����_5W�2h�����v�Km.�ʍ��mgԥc>�UoU�˹5/w}U�6��N{�f�3�d��sc����w8��qg�vN�^T{�>F�?g6��"�TN��&��_;��-��{��Z����3_C8ȟtH���37=��8c�yd&���=I�Tf��dL��;�^��o��,m����\VM����ռ��An��[�� �&;W�#���JM��j"�ֳ51dTA��z3��H=����3��`��|����z��}[��N�uA�18:�I``�$wg�M�6������U���cɢw(�-��Y�qn꽉�/yJ髚�s�O�=o)� ��Ӹ�.��C�\���,f�����:�h��A��1P�K�TN�|�DVU`�=L��p���3���K[�]Ϥ�y�z��ې�����..#U�۬;@��i3	���sy�J�/.�Y���Gk����2��])b���"}�6"���+���N����E���}/CIe�,8��s5qG�L��
�k�$F��b]����d����ȳ�5��ǵC���ۀ$�H�b�$6{���.�zu��b�;�0m&������ˢ��e�Y��`��+C���wX�4Y��<�M���#PS5��TSE�ZC�8���b^,gC�|9̘-��-�6-}H�D��vw��t��z�I|�n�][]}d�ϟ|__}��)�����!/�4{��	f�l1E�ojڅ��Ԣ��f��Ӌ��q;��Jś�����|�x���:D��%��7N��d��]���Hs4構��=��/�+�<)<s��$�V�/����ҎN(�
L՗�b�G9B��y琱M
�TA��#�^������g�Zm�T� �E���}��[��{\�Y|�k4�{�.�v���Ej:�ʏ?n��kQrt���ɧ�h���t���v�Nx�s���y��/1���k�6�+9��~k��ͬ펏ݦ�u�Ϊ�&�-copk�p�%�vޡdM\k�*�e���杧�u��]��m�7:ݶ�N0�^+S�����!K��t�?]+E�a�����S�ޙ���\��_P�dT�:Nr�p�}G6���N5@��s�OX��#8q&�8�<ŗ=���B�_��z�z���^�8�.p}��fhdS���?� �d�67��L�<��Zr�s�ӯR=OH�řX~u\3jӏ�s1\���� �&�q.	� �{Ʋ��g�q��v�ν[ga�޽_{</EIĩ%�R|&YAb%�qJj�����J5���~B;ur�S�I�!4�VP=��iy���QC4����9]ΡQDJb��&�ڮ�$��áX�n��w�կK�=����ε#B.^C v:�[�ץ)���ڸӸ��[��M���ݓ��V�eoaV�˫'�\ߎ�������1`�$�ۊ�۠�^"���v�'{����}����Gv<��rxg���t��8R�����`�l���/<��zbo��xn�!����zr�^"������=�J�#]^ةݹ\�gć���H�-���ܔx�V�/�\��e����h��Y�֙E�<-�	�MO*�Г�{Vr>�]�Hf�LI�\7�=��7����=����E�	�o���e6f��m-�d�W~"w�جp��')���tjt<��z
���N�ш0��>���l;�̤��Gz
�7��q����{OV��<�,�#N����_�(-��{�U�e���K�]w5ЌL��|n�*n/L5�N%�-����[s`�k��ؓuw�M!q�8�/�s�Zڂ�#Nz��qh�
���sd�JtKh�4����2fo���;��N�	Һ������q�G�����u��>sJ&�V�>�Q]��k�i��j5�ٍtne�蝘F0랺G�A]��om�����IG;.��=כ�kK@��؊�[�y���9)浮�j�����wJ�ˡ�Ԕ�c:2f��홭+��z��'�=����L�pq�BqNf:�������J�΋`ﶸ^U�b����3���������z�r1�SE0oU�7�����W��wةe�7�ú��ߍ��O�d��~�렭/[<T�"�Q�j}N�qwJ��>����m���M�`���{��ޓf�����c0F���Z�Z��'A6m⚲8�R93��#�m)8�'ļ:�ť��K�"�n0�D$DRԴ$G*�"��Eڗ#�d��#�>ځ����1�q:#��T��"k)��KO���VJ���kV���G��R��J����c�$f��uFY��1��[�,8C��"=ޝu��viT�X�R�/y���%]m#&oo4YE6���7���ip�`�|j�]�sRxv��Ϫ�>��5�գY��g���z}ϕ�����}�A�绯NΚg�P�{]]�B�,^��B�1��Ȟ���4�n��鳴���a��iO���l	��G���g)�5b�D-\W4��=k��~��MPܮ��Z�2I���r\W����������W{'.�{;|(��a�@�4ش���QC������f����i��n��3��{/o�dir��}��ڂ���e��G��BI�������p�_F���ܺ�I���oo�AL���AFm�<��LqJ��.^�#oU`���Ĳk��5l��B]�������	2���jfw���:�ݦzR{WA��u�Gi����ڵ-��ĤW � ��K5�F:�lU�뷭��m�����s0��܆磝��N$嫈����<�{uܧ-���A�u��h`���Ƚ���H	ٌ˱�s��mj�F5�:�^x��z;g�����zz�U��d֍��۵c�[���$Q	=���>�����;y�^;��z2l�g�	�p��]�/[Lb��`����޹�Yذ3��|��ș����p�Ҵ���ׯh��3�ڻ��OtP�S34G�R��$���s��a��[!M] Ac��Z6�<���,�7��YvS`�L�casDp�m��"x�U�f��݋4-I�����	!��;�Bk�8Q��g��v�ĀH����y���h �����,��I;�Wuco�12�:^AHS7��1�Y H�q9�g�{p��7�hnj%���x-�oUZS�0�3{%u��o,�������*���]����t#��@M�pC�����9��9>0�RUSB�ꗚ��;�a��捁'�����������qd
s�.
.v�@RM}�����z-zf~;���=�s(E+�����~~x�x< ��pL��9� �l}?~���|�l�߽���޳���U�p�r4����D�~}��qy�m��+X��pt���ڲ��P��9&u.Hb��kp̐W(�����s6 [z��w��v��Xʛ����H���@��=�[3��4�.��0�4�Y7��oiї�[��=�<<�2R�r=li);ӳu>C��1�l��H
�!��N�5��n.�ϳJ͏c�֗*�6�Uu�*`o������R3�3o��7d�c���R9�����uN�&��Z3->u�lW��M�Bbh	:,k6m۶�R�Y[���T����Ź��l(g;XN�}C>��Z���Q)�s&�7JkG1vZ���A���\ҷ��|:^�	y3FK`��/a`�7���H��#S/�O���7���N�JX���Lq̼�T�	�=�������1^���&���7a
uӕk�rML�ݓ�� N�_y�\V[;v�,(W*�;׎�%AKv���I
;�v���0���.�o�yrI4d+޻ߟf�?�ݚ�.�z�mGq�^iz@R��K^w�c�~~�/��9f�O��x6oG��V/��	TU���R"�1��ˮ�t0*������S��!�����w9xO"n<-��4�=�65���.i��r\�Jl9�͡O����$Km6|� Yzo���jo��G�QҀ�i��@�/=��r�]�$j!���Y�:zwN_*�Z;�1��a��Ň��o0$��gJ�͞[1�A�z�=:��;z�=���l���;1;-ުU�����to�����ʠW����ue�<���u4Tcv�a�;�8�=sWY�!���A�Np��N�d�`������N�!P)=�/:#� M�,�q��N�f㔸g;��\���e�����bx.�$vg+�&v�lvܛ�6���m�w�߿>�����ǏE�[U���slH��'�$�ϓE�*��HZq�	���
D^��������wOz��޵V��ن������5յd1g�N\ �VK�k'�@�x?(�NȘL��S�D�g&���KV�Z��k�vSg���P�5��2�4�P��nIC� �X\�]�����^�I`�
�8i��6VE%�3H��7����tӫГ�x�k�W��H�Q2R���b�P�I"y3n�<'�y�6<5���LK�R�E�ЬJ����C`���	�'�n!j��_MX8�YOs����apgc̏9���p]�����߉R�ԁȆ����Kt�t��ݘ�H�2J%���-|�L��Z[���'R���ϸ�G�%��A���c��oj妶_Y��=�|N���B��@��Wrw`�6�
�,�6�6���OhV�"''Jf1�SUE�?���ζCv,�,DN�Gm�.�Ȣ�kt��aV3	_�ذ��"���r��tѺ�+�:NZ�Iq�v�z~ɸ&u^�i��J�h���l���%x�?Wz���i|��غ$ጉ�m`<s�`�NgR4�m��s�+B�,c��D$�����L�@�6욮�?�w7���` %�:� 2�` �����iN�s�T��<���x'8�Vg-��K	<O�^L����O�]���һ��m�܅�u3�l��L��׾���I����ڱ�L�qZDip79����~r~_]�����l�j ��e�8�f�`�p��rl2!�l�IO����ȭ��w�h8�?��<�k�}�w���J��H�Hn�xs�Y	c���F�6�Ɲ퐑���,L�#C_I��p���h��})�X�ܦ�Nm��ps�J՗�*h�mgw9�hq�y]��d�~��a�!��KV����u�,]��&ɩsh'����o�F2RG����=kNv�E]�zu���7M�ѦS��o+�N�LjnL��lMl�9���w[�󀈢$����Y4�9�=xy�[��i7�h�끊2bp�j�R�{i+FD�hV�fT��<quu�%�Yo{�[���:���MɞJ�V��K�9#k�;���wǝ���v��ղfsLM����������hk�F J�)yW�7^�v��#;Ѝ�fH�Z�Qz)��=ph�����S�`΀�W�LX-J��t�3v>��O���y��m̖-�YԆ��S����^���v_��3�6k��1c�첟���J���(�TҷNv���#���AvZ%J����:��qV���wGV�"��\ Ýܚ��ח�+Vyoj3�+���_"�j�k�V�����g�����[��K�{sHxޯ
�8�O�X�yc|�ݝ!�Ⱦ��lw��OO
:at"���l}�6�+�P����t"6+����xr�+j���Q��\t��t������,�������/f�b�����I��7���=zxo�3zp9�:yu��h��(,���з4PМՐf�/�걊��e+�z��p`��.;�X��ޗ���ϻޗf��ڳܤz���`Ȧ�R���#�R�M���oߥ�t���R�v������T�7��y�V��ϭؘ3�Y��s8��}KJ-�齁��d�� ���5_�I$�J�����FKv����s�i��lə���\������fֆM��5���on�a�;n��naT����D��Jը��(gp�c��uu�=r�ç���6m�T3��^�rg+��<��7+���<�����-��V@��ĥ��yK;y���G'ϛ�|7��y_����\�\r�c`}8�e�!��F�J�Xݕ<�p)X��MN�3�2�=�V�;�Ա�Fz�:y-�w0�W�]1�,<s�zݥ��w1��;�f�Cie�m�x��WF�p���<:��wK�<���<��.9���qn̝�W�ٻ"ͼ���&��n7ff#r۠��ۇ,��yy몼�����糀�&+��h#�öM>���Y�Dq��>�[g[�F��v�Ky��q�q�k��܊��͸��y�Ʌ�N�	��m��3Lj�ё��\V�e��n8X��ݧ���m�8I�Mפ�1�����X�]g�R񬭸@]+�sr=�y��}���a�8�k6��]�&;SskS:c���q�S�g:,�C�&s�G����q�O����w����_��ug�A�`[on��Ƅ�lk�ܝ�ў#�ۧ&ͦnz;F�{8��S� �q������C�֎�r�q�\�՞t���`��u�[<���GY�c��q�<lloC�J���S�&��u�^nݬ �C��i-����Z� �2voW�+����K�����H0�Ӱ�}�gn���0�D���U��{����dP��X�7dcCg
���W��(/dm�^���G�g=/̬���||9�Ԏ��Q�vou����}�=7�R��Ǭ�+�2�\��R��ÆL�W-��U��L�e'oX�b�ŝ_g��h�֒\�2�ݫ~�g�����g��,�KQHv�ԹW7lܯ=U�'��|��@�Yށ�]�Ц�(�x�j7gp��OQ�z����L]w�7d��H,Ⱥe��h��2R{���r�e;r�KW���k:��o����3x�_m��jĆ�{��ۼ{_:XU�A�" �Go����3�g_
Z��Ѵ�7���Nq(���Q��Rr��5gƛ��s�-�o62�`к��(4��Ԥ��c>Z���Aްe���S yJ�$�Y�K�"�w&1̭�YW�rRw� �
?7Nñ+�Zu�{[g]�>:���P-�%s�+��=�����"X��ʏ^&�|���Kz1ȕ����y��6E�J��(�;e�VGFe]��n���W6[<c_,[�Ho�I�hqo}8�7�ت{���j[Uon.�U�����=!��۲B��e��v�]��b���N�����0��͌.�����ݺO7���	��M�.��sve<�.�Q�Qٕ�Ƒ�l_B�&vv�����!{�GC�l0�ҫ����!����뺖�.ނYR�9�H�ʹv-'�f@B��e�pT��Y��`S�猆�gƻ%�y=�Lܴ:a�#܂�L�u1��[��#�#���4��^&X(����u�y_��W�r��7�J�r�7ј�Y�O�)���Bg��n�P�퇈7I����B�㵴i�#�2�"�1m'�Nηt�"��qїc��;E���oM�z�H�5�g�^)�l��xy�_o��Mev#.�E�9���.��)�h���A�y^7TC�����s�:��Y�}t�ڔ��Z
8�ۏZۋct����V�w9y���fD�d�H����&s��Jg&�1�F��.yfHsӭ8�_�Uj��a}�o����c�*�.���̫A���
5ëi��=����s|u?D)IgbMa9F]�D�!�5gF�]�w��vI���+/N�'��t���i�6Yk.8{�=��K���H��8=��f��&m�7�ו��$J;����#-��N_u�b��N����~о{�����N���3t��0k� Z�ݾ�4w�����a��ӝ�qk�Iы��r�����\��. ��e琜i����/Lm�-�����e�[n#�q垺1\���on3����2�W76���٢i�b8�"��rk����^67n�8�,�k�DV�U�&��|�i�s���ֺ�}`ގ��EP�u��P�؇6p�)'�!�k�ڼ�3�;�iXB��V��r�xE�<� ���@�HX�,6�DZ��[���9s���4/�H���4t��������O��g�p�p�3���]�~��Y@Rl-�"��,�k�M`�פ(&DS>8���zq3�fl>�����T�M�O�bά�5/��6�[,}��1�MÍ[�/f����sj�咜�ϓL��1W���=� ������/|n1wI�$B�[�c�pI$o>����������BYbڴ���q��v��O��j0�k鷇98��s:�;��{6N�e��;/�]aId��mV�}�P�g8֫�W>�1����
WZ��#V�B'��ڵ�~��������=��L�IE�p��10�;�tq�Y�O�\	n&�}�E�=�&�tt��F�^�)�Po����Z�|��<������%�L!�W��{�(fx��Q|zr�4��sF#�d5z?����-9��}�lܜ�5�s\Bvp��7j+�	[9�f���'b:�b��r�k�O.��u�+	]c�:OcA&�"D�{�l[��4���Q��fǦ$"u�	W��!���--шk��8Л���7�m�O,Iz#N������X��Yr��G�k�N"�n��:%\+5r��x~���0y���Dt3������nq���b|��h��F������"�
�8��i��X��ݫ�l��\ۉiష�����T<�B}��q��.\8�"=��,�Пu��z���0�aQ�L�*�#j�g��[�Hc���,`�wZ#O>�c:Su�ť�$�9k;��Z�n�W��+�c:RY~E,������pM�t��ć��a#+�fx�L���/n�~����r�+�J^���oJk���C坩B1��;�:�&%]}����Ph�dt�T�2�5	��!����[V��ec�^؆�guN{��o]jJ�s����3R�r��^3G����l��&�n�g����َJ
M�^�>���d�ŏo����>���w� ���8�����ޘ8n��/��7xWE��-���\bk�/7w��*J&�Ű>X�Ʊ��5i�2L-TR�4h�,��AR>�_Lћ�m"VV��9$�]6uu�q̌�;	VE�HJuˈ�Mk8�LID�A))��`��PE|f�j�UR��1���XUy�CꑥgN'�}�&���Y�H��8�A�3�_K��&�]Z�?+|Tj~��]��Q���o�u�������(T`��kUE�;U+�Sk^u����o�i�����>��>#�,:�mm�v�eͭĴ�[�wk�벑���:�|�)�h7����bsԛ��U��g[vu�m�a�:�u�G����۟�oTە��u{b����i+�Ml�x�s��wW�W>���s��AE�7MX0L1�� )��fg��iO7��H6���n��g99I��["9�!��UK\��HR14�a��u�߿`��y�����k={'�����ʩ��u��Ã}�49 �z�X���G�^��k/ha�pr@�>��iMb��;j�%��\�d���Q���_�ٷ]9�QC�N"�r���J�âq% �<�y&uf�\FIod��N�A�Oʵ�=��p\�]�vf���~}�~��M�ۑ�tu����5�=�ͮ.z߯���|�@U���cd
���ӿ�}e�v鍮�z��f=i����-F��㽗v�r�4�8y��{|�*=��2v�]��F�Qށ�2��γ�r���̯�'^�2�.k��=(6���/��KM4ϸ�y'4�y+L�>��~�{}��}�a:�)���̦�XH>贔���s��sْ�g�>{;���f"���+�=��մt>l��M)��4�;}�R
�����Q �[�ƚ�c1�D�I�Yy��S'�Jk��BH����`5�%��iɸ{\�P�u�L�bC��>=�op��0��d�1��m�E�`<W7&5�d=��k�C����K��j��;�\��\��v ,M�����)�MiJ�,���SZ���}�Y����=���7���CQ�M�����`kq�.D��e9OS�3��NHj�zV�0�/�W7*Қ���c����bZB�`*��9Q8����-�5��S�H};6����ΉE�N�����0ە:gI�N�[߮nfM];:�q��
�p7o���3�vh3 �f��)cc��f)r�p�FFZɚ9��8yk;r��!�b�Vs̘�ug)Xs��/Z!��x�5��׽6�C��Fh��HU���a��&q��U�u	{����aB�ҫ��o�8q�w_��&v���L۪�ݨ�u���T�6��pIrw��'��P�P�9��y�oR��V�sv^:�N�a�-+�2�����$w׆lؒ�·r���$L���+B�|����+�w��8#|���Aл']����U{�wsT+x���ПY�6k��˪M:�s�sh[bu�3Օx<��{c��]n)���f���GOLGo�x�{��;��&��\E�U�Af0�eLp��H�����CM#������i�-w0�R��V��ޓ;�`���A���;�W92�uɗy0VR%}b+��u��ݳ���8�w�-��"�,�h>���k:�m�;�����ry�'���8,A}�Lo��o\�=�☼�΂'&7���8;��H�2�]�0���N:���N\0���F/�� `�@��l�ec���%H<���2��񮴓
Rb������L����*�X��PjX��[��a�ףb9f���]Λ��Iۺ߯E��Z��^�Z��$nb�'Mg����[n���9..�7$�����`	fݯxq
G�@��7��|�b؊}'�
#vz���u@�'7���Ǩb���f��m-��+=�G�@�0#��__$t*+��!�!(H$#u��CHz �;�]�]���ɚ|���1�6� v�8Z���PG���'���}��U�� ��ɚ�f<�w�eh���/�f�/nBܐ1�է����F���c��|�<��b�N��H�N���^�� b�WU�yL:�"(��\�)icc��TY�C��;unL캥y�-3��2��ލpz������{u{K|;Dt��8{V�ݚ�����*�W]��8��w[�H���'���ɶ���<�^��k�W�[��秱ѝ��-IЈZ��uQδ�Po93��Nⶴ�/�Lov$6�ײ%XH��/�:�c��y�����^���Ajv�%��PS�.��6����S${q�	��WO�����)��ȁ���+ٔ�6�����*��o�)A�K�����Ñ��h���oy�b��ﻠx}������kL-�V �|CxM�A1�gR�,y��qkb�����$ձ1'.����S��2��]}�\�XV�7��<�B�g&k���ϒHUwH��<+6���{�p�<r�g�a!�Z8�G1�4:@�u�4����L�vݵѱ�+�W�z���#O�<��#���'�~�ghm��^;E�5��Ö"���B��2��@��Q��@���Owd�U���TJ�wrYu�
1Q�;Wp9t��az�ggi����n�G՚;ނmއ���V��\�d1̱��l�[�u��ƣ���J�r�%�O
:Y����9�w")F^�ni�%�٥S��.Uw��lÝ�E��waYj!jY��}����P7m�,jw�"����d2�Q{ x��iOw��UWW �"�l�ϩ
ׁu!�ۍ�LB���
�ˌ�kb�테l��ǈ��h;u	�^����	h�AZ�c*�>g���YJ�w�����}�	�a7�k1�F�b��à�� ��(nn���.*>��OKȶ����$���u�Toʁ,�Wqdl�$�ݛ�ۙv=�O�ToHv�G����ޱ/Rg\ַƌ��]⮥��=3���2�:1�z��ڱ��(���I,]�{2��c�Fu�%gg
�;m����sZ�sR��j�ˇ�P�@�O�\���f��:3���#��;w��ҩ	��n�Z������QdMƣ���NLfˡѯ�� e4]�[ij]J�hwp=+�B;��<�-�h񱎲�� �J�i2p���z/m�ڱ��;��Bi>��a�mX���93;�>�b5D6����|��R�oqpu��g�`�c��� ��j�wR(�-}����xt�t�q���R9�:��-ƞ�O'p�{�^�TA4��R
�Y\�� �w5jf�V"���Qx�m���TFr�=s�x��2��S�';W}>я��a�{
�������jx���[u�2یK�Ce40�	��Q�ѪWqsޮѬ*�7�P�{f�Y��j�hh���#�_m�3�w��^q��;�@�5;�m���n:�G��Vt#�{`�Bt��"qM�Ed��W��Z�Y	!b�3v�[{�+����k�T6���WmĢ������8��<�L�\����(8r�f�b=��.B�d]#�8��� ��sJ���㋀�p�y¾�c j��^�����_ODm���е���}7�������}�xB�ɤ���䵙"�}��K���ݜ���zm���=��*5��Wx�;�X��Z�<6��=m��8��3���zwf���,���x��v|��]�ݫt�]o�j';tڶ�l�Tw�b�c����sə�<
�����iٗR1<]n �!��3�`����zUI@N�c8���n7޻nʀū�6������6��Ed'��޴tSlk�`�zKDNC5�h;x˷��ܖ{|�ǉ��{���ޏ��ٍ0M<��$�fm�Uq{%������i1��l�sq�ݶ{��X�^�.�Y���},��!u=9��`͗@~e7����'�-d��#H��1��Q���;l����Ϧ ���]# 3Kgg8N6��q���ݏ '��0R�kO��,�OP{��*�G6x�މ�����i�Ӳ�Bڍ�#J���_�nh4���u>��3�����y�خ�gwu�o+�ø��we��
m^�>��W/���v�K{m�ip_5��L��޵� �^l?r �G��;cڇ��^�f�֔(]�.�WG$4��ȕĪ��>�]�xR�BQ��,,��a�7��z�B���vn��A����Ίx��ݔE8���U2��F:�u�>���G�I�M ��^��NN�&�'\=T�i� �璘y��L�ݦ�L�	�C�C#�B�[x���0�[-�uM�����7��vy�{�Bo�l���K-{�O#;ۏ�qe�GS8
���矆I�ױ���.�8v]��4��>�h�nv�<A�Dh�+U�s;�pg7,-����ʣC1��P��*�+En:�h`�"J��K�5�!g��z7rՅkYmt�Y�b���v`/v������~4��9���}��H����F.̡Y�J�&�OV���������gsڹR�g5J�q����WV/�g����N�|� �L��f	'N��
9����u񼧘;L���"X��Uo���F3@]�7�@\/OK�\�[@g295\�<��-��%�kx|��g��G�����b�,����0�K
���e�{�/�,HA�؈=4p��h�H�Ƞ	D�b�T4��ل�$۲���6n�h���&���w}=�������S-o�B���6��!�zK��c�N4`�M�F�wK���*���QQ4�Am���w��������q!֞�.�o���ût�-җXh,}�����B�Q�������P=ޘ��V%�JP�fGq���8<W�]����Y٪i^���h��pV�Ęo���=7
D�W�֣)}j�Uic���zo�*jkh�E�;�:��J�8����<'�v��3���3���z��C�Bt{Q��1������[Ȝ���)Mv
�\YxZ�5s*��|��nj�y���=Ga��s��@���!$	$��aB�����z
 ��9[C���c=�]T7:�x&���AQ ���Z���@��l�V腐֯X̸o+w{\@�&�P$����.��ʪ$P$ I��!QV�
��7"U�Y��(�� 
�*(TUDd�f�QV>��#J9��)��m5���d�:Q�Gs݌q�(2@12�@�/������d@ D!��t���W�
�����&������nv�Z��:L-?��#]}������c8��n��?.ރ)G�;�/y��t���?�����=�D��m2�Ҟi��&�|��aObw��ju��ǣ��0yn����
  v�ܴ����;������>�O�Q@@�@�W@�)`{Ǩ�������Ѱ��Qsg�?��?���;��� ��t���Hkνp= ��
  y���D�u!�<��������@a�i�<� v6��v�"�oN8Z@�C�o�:��`�*#�Q��_��S&Dl`ِ1w�D�|JP���-N�Ń�Qيf���ǲ)'�>S&��9���qA'Y/�PT@,i���r��}"� [�b�D\QHD Q��X+QA`�i�d-% ^/bB��v��z�p��(�������h�S��t8����!H����4R��!�P��/��� x�t��vS���6�H����z��u&�û�/Z`�o�t8<��4?xp���+���Cԟj'��������C���B
���}qp$~��0��pN�O�^������}�I��7�ؤ��,�]�Qk���N	���=~�>��u`�i��e~3��$��X1{����P�7> �|}Q�=����K�z!0�4���O�z�>�k8�{�6I͛���J�s�"��"�,�� � �a�
  �X`>e����D#=a�H4l���+��'�rᬥ��d�aB��2E�0�ꔥPR�F@�?�d�Hy��}_��׉M����^)-HhMj�~A�9��p.����o������B��P�+��G�3�����B�:�pF����Z������l�¹401A��+ � ]P���'�n�=܇x��
  {���	���r�w)�}a����=��z���2~����77���Z>��>c��[p:`%)A����}A�I/ʿXu�5 ��KM��	0���`��xl
  ci�;?"A��Ċ>��A<V�Q��pȟ9�(�c�:������U����>�1�S`;�	��O��o�k�h�҅$!G�������T����w�tt|��s�=�}�������x��K�dO��.y�㳯����q��ĩ(�_g�z;Dɩ䧙N�Y��EɃGYܐh����;'��n���`{^�.�g��k�$d�s�~"}R�6�z�'�У�h0��Ά8�w`�S��z��@@��P�~	�ꇼ{���Y��e�HY	�p�t��8P(�8y׸�l\'�=!j^�'dP/�S� ��C�x���;BEK�@�j$!�w�!��.�p� h=�