BZh91AY&SY���� �_�Ryg���������� � �
?|�/�ݺ�Aq�k�    �4���dd���0�4ɀi�4�ɄM a4i� 	MS�OR��4i�ƚ #&  b0"T�zOQ���4��� �   2�&j�jz�4�4=A��@ h�M �"ɠ!�e7�S�i<��=L�A����PtbD�IG��Q-"?��y]�H1$��1�8w�H4P���&ͯ������Z��BWKm~��� �t� ���f�@I�3IIT�:N��:j8T6+M�kP�ѦUhc5͔�7j��JT���R2���W��%V�-.�󽟺���v��3)%ԁeZ@T�wo��g��mRy���e��EбU�M��m���V諒�K3@)�J}�(�E��^߆f]\�l����x�\6����nAP��L��!�����EW	Y:%q�Ru�o��
���n�;1���[T�0,�]�&	�e_������zjt�-�n�ڇDq�2"��R()�
ĒA��� �,I$�i�v�5Mc)��&�ӁMu������_� `ƈv汭կV@+x�m��n���p��(Y�{���eCD�R���,�i��쮫�`֥�М�ȥ4����+&/������Р�ԍ��[5^M)�1Cm�u�kK��y�9�՘Rb�ε(���ݪ�g3}�8^�e��(�M,��r�΢��C#D�|4����*C5��N2�~6Ҫ��{P��*5��A��62�M�m��`۪|�R�R����O�{R�UI�E6y��`΅�W��IkE��ɰՋ61def_��kg�x/4��״KݍeSZ��f&V���/6uX`|mUi�~�J��ZN�{��C��Vf�l\fVe�*�*�B&���ZF�'�J�d�Q	&�؋�CJ��H���E�G&�ɘNE��"BPU���I�^ȏ8���@¤��Q����Ј�+�@��������g#g��
Lm���[����Z6Y�e�N.eZ�<ʥ=����ɒ��as�{'b��zu;e���x��R��cN�Q��G��M�M��I����|��M��$���!d.<#���>������ �u��<e�;jw��?#^���.�ֽ���m�?Gg�3����oU�甾'��+��إ*9���%����*L6�>�*�u��lCf�b�^��	���2G�X�qR�/I:BjRBR����gM"�M;]��s��o�з*��`��A�)�3����T	fb&�ԸSC�d�-/YD��b��E(2�e�Z1��̢��׌|�����0>�nؼyuF��ԴeP��R�-Q~nXg��ȧ6�ɤ-�z>�I����S�cq����*�/f����/0C���gӼa��>s�C���V:C��%�0�;9�&�EF1;�5��1�����N�YJ��fqx�)~�����;%�2#��]M�.�Mݳ�35��OSk)���Tl�w����]w	��:Sg�ɳ]UnN�~���U)�����T���3����s���mO��'c¦R�)R]n�]�������TvE{���yT����#���C��5)�H�G!��w�&Q:�E�Z����R��\��ޥШ�_����-$K5CL�<����H�=-O�d�Ք�}�ƥ4�j0T�V*�D�6���>ׯX��dl�D��Ȥ�ZM$��\�j���ֺѱkl�*ee�E�6,aQ�Y#	QP��=��[�='���J�8Ga�q�l�<c��z���{gT^�68}�}�y�g��>�/��o͛�D����G�K��^'v����N�B�[t��>��I��t~�+�&o~�U���5XG�ss�8�:1����.a�o�}����ĉX��%얔��q�RT�!q�"���6���%OLj��^�S�KL�N�IS�� ����-cJ��*K{{{��3��xek�z����v;��8�#û���7)�Z6dG)f��Fwd���3�+�b�*����%qߨl��Y�㢨ʕ��Y�I�E�	�R�sj�M�/՛��j�1�&ݮ�Yi8��8���h��fI9/�赹{��1��9uRJI��"��0�z0G\�*H�R��~���L�)<]N��94��c��0��QƊ��_�x+�l�?/��ǿ�d�4�P��� ƒ2�����'���)���