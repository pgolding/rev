BZh91AY&SYç� ߉Ryg���������� � ��2���G}, {�B�wq�v:��@m�� ʅ�"��S�)�5�&����OP���� M0d�52A�# �`� ��1 h�Sjz��ɠ 4b   HD ���zJi��Sh�OHb  �RBz*~��g�yO���C�@h@  ��Цh�S���hb��ݻ��H�ڈ�?�BY~����"�2������Ot�WT�H@X��?6V�-=�?�t�l1��D!s�U`�|��[q@Hm#�?D�g0����zT浲��GIt6JJURGUCN�Hj��d!:�P�Ad�ʙ�Rp�u��٦4&i&���}��Vf`ط��e��#�aL^[E��bTI%�b"������	���qp7��^��V��\���@� #1)�Sv
lA�L�]�0�Ƌ6���j:=�G����Q�gL(���)��!	���=pƵmFL�Y�#B!H�{O�ȟ�ܞ9wޞ�׼t<�2�F �]�J������Ϭ�ٱ�nA�,0פ���3E��1�}|�v�����(�U�=����<�zs��"-C,7�(���G0�b��+�VWgk[;I�G��ZbD2�����a[r""K%-��+n���WI��X#)Z��Й�cLj��'�1����|}��R6���m\
pR�V�u~���υ�xr�5�)#b=R|O��G�@��XuFd&��9�zq��
y�1���'��p�f��4�8�dl��������j-�sY�xk����[AnՀ�8n��d}8�RcDxcËf\怷��GjA�6�M��C�]�iuc���a��d�]��:��-6��R<��]x�/���.���@at�gl��bu�crTaƩ:�η�ŶJ���y1K|�w�n�h��5����m�.�s1��c�N��3`΋��vcP0�ngTL=��(���(�t��vW�h�N��(�%<#��$B"�'\�X袍�["��!��+���fCc2�47i��m�m��$2	1h���y�5K�ޥ���T�ʒ�k��b#c�m�ll�@t�YL}�E��cKvA�h(�1��3U֬���Y@���s7Q�z#b�5F���9���AX_6�����$(��g��M��K����Crd��8�"�b+ h�4#c1,����GH� e� �mclƋے�mu�_�����q��m��^�Y�G��R����0�����9ѺN��#���
,�Z����Jh-��N�("EGB��HFZ�$������*-
�$�S騻
a��ݑT������R��3*����M����!�����c�aH�<���ثU�.(x�}7diQ�ȶ�x��T����_p?�_}^��"VB�)	�`T�����6M�t|<T���;"t쐽�5�.�����i�kur�՚S����m �@b�e�L����5ٌ
�� TW�K�+��<�/e�}k�U]��c���p��IJ�Q�k������א����.I7tU.����ѪHժIVv俨��hLnȐת������ ��U/�/���̏�Z���󜾺�N�h��d"�-�`A+��?g�qj�=�x��݀4pZ��$a*��2����!�7c�FQR8,�#&4�H�E&@2`ab�p�_F��{K(���U[f�*�ǳ�qf��h¢UIU�9V#��4�&�R�6�D-��>RE�>\b�8��EMݏ���)���TK��.7��i�:tƔ��ˇD���g˞��=�o�O,Mb��( ���:�щ%�){ՠf���6O'�����)��C�s8�[ڲ�$�W�k����B�8��E"��e � ؇}�-N��2�;��i>��۾N��N֋������F ��6������S�!�$ќ�qB!�51�2 ���7��7y�5�P���ꐤ;�3��(�*\W��k"J�W=����$Q�OK)T�Y뵈���E�U�wɹ|I�5N�C�ah�x�!��Dy&)1��_��J������*UJ%%I��^(��,�t;����3�=�EȔ�4g��0��$�;cH����Rl4���ilKL��
j��2�"!��K���l,Pt]h��ֶ��`�I�.���aT�'��E rn��\: �H8 [I�)��Hz�im4����uX�޸��X-���ɔC�>i�Z8�I��wNB�H5�>6�@�렘��@�9R���[����c�鋹��&�������;�
����4���ұ|Y#�#�n�����gզTRi�7�{*����d�:/>F��u*�B�j��h��*�C�:QJ��]B�-hX�$��wXaQ��v�dK��~G%�����d��%O,��{g]�˻O�WFe��b���Àzͺ��Τ��L`�Zy�>g���9�*Պ��.���/V�i��_\�x���)��5ԇ�N?O�t��Ո�5C�-Z=f��Ŕn�a<P�m�?�������yxl ��a�at������FT���M��%�~�%2�����wf�w5�Oص��\�Ք��O�#��wm�f�{\��4/�&���0��i����0ݾ��z5@�ld��AB>���"�|a�o�:�6�I'YE��d��eM_::DY�✇)�1����������]Xj$��$��G���������.N#L��K 0h`.&$�a��`��)�8�8